`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07.12.2023 16:07:01
// Design me: 00
// Module Name: instruction_memory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module instruction_memory (
	input  			clk_i,
	input  			reset_i,
	input  [31:0]	iaddr_i,
	input  			ird_i,
    output accept,
	output [31:0]	irdata_o
);
    assign accept = 1;
	reg [31:0] data; 
	always @*
		case (iaddr_i[31:2])
		                                          //32'h      MachineCode  ;  //	BasicCode	     ====    OriginalCode

                                                  30'd	0	: data = 32'h	00000013	;    //	addi x0 x0 0	  ====    	nopamoswap.w x3, x5, (x1)  // Atomic swap the value in x5 with the value in memory at address in x1, store the previous value in x3
                                                  30'd    1    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2    : data = 32'h    00000013    ;   //    addi x0 x0 0      ====        nop
                                                  30'd    3    : data = 32'h    000100B7    ;    //    lui x1 16      ====        lui x1, 0x00010
                                                  30'd    4    : data = 32'h    40008093    ;    //    addi x1 x1 1024      ====        addi x1, x1, 1024
                                                  30'd    5    : data = 32'h    22222137    ;    //    lui x2 139810      ====        lui x2, 0x22222
                                                  30'd    6    : data = 32'h    0020A223    ;    //    sw x2 4(x1)      ====        sw x2, 4(x1)
                                                  30'd    7    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    8    : data = 32'h    333331B7    ;    //    lui x3 209715      ====        lui x3, 0x33333
                                                  30'd    9    : data = 32'h    0030A223    ;    //    sw x3 4(x1)      ====        sw x3, 4(x1)
                                                  30'd    10    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    11    : data = 32'h    44444237    ;    //    lui x4 279620      ====        lui x4, 0x44444
                                                  30'd    12    : data = 32'h    0040A223    ;    //    sw x4 4(x1)      ====        sw x4, 4(x1)
                                                  30'd    13    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    14    : data = 32'h    555552B7    ;    //    lui x5 349525      ====        lui x5, 0x55555
                                                  30'd    15    : data = 32'h    0050A223    ;    //    sw x5 4(x1)      ====        sw x5, 4(x1)
                                                  30'd    16    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    17    : data = 32'h    66666337    ;    //    lui x6 419430      ====        lui x6, 0x66666
                                                  30'd    18    : data = 32'h    0060A223    ;    //    sw x6 4(x1)      ====        sw x6, 4(x1)
                                                  30'd    19    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    20    : data = 32'h    777773B7    ;    //    lui x7 489335      ====        lui x7, 0x77777
                                                  30'd    21    : data = 32'h    0070A223    ;    //    sw x7 4(x1)      ====        sw x7, 4(x1)
                                                  30'd    22    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    23    : data = 32'h    88888437    ;    //    lui x8 559240      ====        lui x8, 0x88888
                                                  30'd    24    : data = 32'h    0080A223    ;    //    sw x8 4(x1)      ====        sw x8, 4(x1)
                                                  30'd    25    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    26    : data = 32'h    999904B7    ;    //    lui x9 629136      ====        lui x9, 0x99990
                                                  30'd    27    : data = 32'h    0090A223    ;    //    sw x9 4(x1)      ====        sw x9, 4(x1)
                                                  30'd    28    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    29    : data = 32'h    000100B7    ;    //    lui x1 16      ====        lui x1, 0x00010
                                                  30'd    30    : data = 32'h    40008093    ;    //    addi x1 x1 1024      ====        addi x1, x1, 1024
                                                  30'd    31    : data = 32'h    0040A503    ;    //    lw x10 4(x1)      ====        lw x10, 4(x1)
                                                  30'd    32    : data = 32'h    30200113    ;    //    csrw
                                                  30'd    33    : data = 32'h    00B02073    ;    //    csrr
                                                  30'd    34    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    35    : data = 32'h    0040A603    ;    //    lw x12 4(x1)      ====        lw x12, 4(x1)
                                                  30'd    36    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    37    : data = 32'h    0040A683    ;    //    lw x13 4(x1)      ====        lw x13, 4(x1)
                                                  30'd    38    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    39    : data = 32'h    0040A703    ;    //    lw x14 4(x1)      ====        lw x14, 4(x1)
                                                  30'd    40    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    41    : data = 32'h    0040A783    ;    //    lw x15 4(x1)      ====        lw x15, 4(x1)
                                                  30'd    42    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    43    : data = 32'h    0040A803    ;    //    lw x16 4(x1)      ====        lw x16, 4(x1)
                                                  30'd    44    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    45    : data = 32'h    0040A883    ;    //    lw x17 4(x1)      ====        lw x17, 4(x1)
                                                  30'd    46    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    47    : data = 32'h    000100B7    ;    //    lui x1 16      ====        lui x1,0x00010
                                                  30'd    48    : data = 32'h    40008093    ;    //    addi x1 x1 1024      ====        addi x1, x1, 1024
                                                  30'd    49    : data = 32'h    04008213    ;    //    addi x4 x1 64      ====        addi x4, x1, 64
                                                  30'd    50    : data = 32'h    0040A023    ;    //    sw x4 0(x1)      ====        sw x4, 0x0(x1)
                                                  30'd    51    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    52    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    53    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    54    : data = 32'h    F9A4E037    ;    //    lui x0 1022542      ====        li x0, 0xf9a4dc93
                                                  30'd    55    : data = 32'h    C9300013    ;    //    addi x0 x0 -877      ====        li x0, 0xf9a4dc93
                                                  30'd    56    : data = 32'h    27DEC0B7    ;    //    lui x1 163308      ====        li x1, 0x27debf5f
                                                  30'd    57    : data = 32'h    F5F08093    ;    //    addi x1 x1 -161      ====        li x1, 0x27debf5f
                                                  30'd    58    : data = 32'h    00F00113    ;    //    addi x2 x0 15      ====        li x2, 0xf
                                                  30'd    59    : data = 32'h    800001B7    ;    //    lui x3 524288      ====        li x3, 0x80000000
                                                  30'd    60    : data = 32'h    00018193    ;    //    addi x3 x3 0      ====        li x3, 0x80000000
                                                  30'd    61    : data = 32'h    F499D2B7    ;    //    lui x5 1001885      ====        li x5, 0xf499cae9
                                                  30'd    62    : data = 32'h    AE928293    ;    //    addi x5 x5 -1303      ====        li x5, 0xf499cae9
                                                  30'd    63    : data = 32'h    5D4DA337    ;    //    lui x6 382170      ====        li x6, 0x5d4da3ca
                                                  30'd    64    : data = 32'h    3CA30313    ;    //    addi x6 x6 970      ====        li x6, 0x5d4da3ca
                                                  30'd    65    : data = 32'h    CD62F3B7    ;    //    lui x7 841263      ====        li x7, 0xcd62ecaa
                                                  30'd    66    : data = 32'h    CAA38393    ;    //    addi x7 x7 -854      ====        li x7, 0xcd62ecaa
                                                  30'd    67    : data = 32'h    F4DD0437    ;    //    lui x8 1002960      ====        li x8, 0xf4dd0029
                                                  30'd    68    : data = 32'h    02940413    ;    //    addi x8 x8 41      ====        li x8, 0xf4dd0029
                                                  30'd    69    : data = 32'h    00C00493    ;    //    addi x9 x0 12      ====        li x9, 0xc
                                                  30'd    70    : data = 32'h    F82F4537    ;    //    lui x10 1016564      ====        li x10, 0xf82f3f90
                                                  30'd    71    : data = 32'h    F9050513    ;    //    addi x10 x10 -112      ====        li x10, 0xf82f3f90
                                                  30'd    72    : data = 32'h    B81585B7    ;    //    lui x11 754008      ====        li x11, 0xb8158480
                                                  30'd    73    : data = 32'h    48058593    ;    //    addi x11 x11 1152      ====        li x11, 0xb8158480
                                                  30'd    74    : data = 32'h    AE889637    ;    //    lui x12 714889      ====        li x12, 0xae88946d
                                                  30'd    75    : data = 32'h    46D60613    ;    //    addi x12 x12 1133      ====        li x12, 0xae88946d
                                                  30'd    76    : data = 32'b    00000010001100010110000010110011    ;    //    DIV x1 x2 x3
                                                  30'd    77    : data = 32'h    00000713    ;    //    addi x14 x0 0      ====        li x14, 0x0
                                                  30'd    78    : data = 32'h    00300793    ;    //    addi x15 x0 3      ====        li x15, 0x3
                                                  30'd    79    : data = 32'h    80000837    ;    //    lui x16 524288      ====        li x16, 0x80000000
                                                  30'd    80    : data = 32'h    00080813    ;    //    addi x16 x16 0      ====        li x16, 0x80000000
                                                  30'd    81    : data = 32'h    00000893    ;    //    addi x17 x0 0      ====        li x17, 0x0
                                                  30'd    82    : data = 32'h    80000937    ;    //    lui x18 524288      ====        li x18, 0x80000000
                                                  30'd    83    : data = 32'h    00090913    ;    //    addi x18 x18 0      ====        li x18, 0x80000000
                                                  30'd    84    : data = 32'h    00B00993    ;    //    addi x19 x0 11      ====        li x19, 0xb
                                                  30'd    85    : data = 32'h    F413DA37    ;    //    lui x20 999741      ====        li x20, 0xf413c908
                                                  30'd    86    : data = 32'h    908A0A13    ;    //    addi x20 x20 -1784      ====        li x20, 0xf413c908
                                                  30'd    87    : data = 32'h    0DFF5AB7    ;    //    lui x21 57333      ====        li x21, 0xdff511b
                                                  30'd    88    : data = 32'h    11BA8A93    ;    //    addi x21 x21 283      ====        li x21, 0xdff511b
                                                  30'd    89    : data = 32'h    00000B13    ;    //    addi x22 x0 0      ====        li x22, 0x0
                                                  30'd    90    : data = 32'h    80000BB7    ;    //    lui x23 524288      ====        li x23, 0x80000000
                                                  30'd    91    : data = 32'h    000B8B93    ;    //    addi x23 x23 0      ====        li x23, 0x80000000
                                                  30'd    92    : data = 32'h    FBCDDC37    ;    //    lui x24 1031389      ====        li x24, 0xfbcdd417
                                                  30'd    93    : data = 32'h    417C0C13    ;    //    addi x24 x24 1047      ====        li x24, 0xfbcdd417
                                                  30'd    94    : data = 32'h    00000C93    ;    //    addi x25 x0 0      ====        li x25, 0x0
                                                  30'd    95    : data = 32'h    91240D37    ;    //    lui x26 594496      ====        li x26, 0x9123f832
                                                  30'd    96    : data = 32'h    832D0D13    ;    //    addi x26 x26 -1998      ====        li x26, 0x9123f832
                                                  30'd    97    : data = 32'h    80000DB7    ;    //    lui x27 524288      ====        li x27, 0x80000000
                                                  30'd    98    : data = 32'h    000D8D93    ;    //    addi x27 x27 0      ====        li x27, 0x80000000
                                                  30'd    99    : data = 32'h    80000E37    ;    //    lui x28 524288      ====        li x28, 0x80000000
                                                  30'd    100    : data = 32'h    000E0E13    ;    //    addi x28 x28 0      ====        li x28, 0x80000000
                                                  30'd    101    : data = 32'h    80000EB7    ;    //    lui x29 524288      ====        li x29, 0x80000000
                                                  30'd    102    : data = 32'h    000E8E93    ;    //    addi x29 x29 0      ====        li x29, 0x80000000
                                                  30'd    103    : data = 32'h    1AD0CFB7    ;    //    lui x31 109836      ====        li x31, 0x1ad0bd45
                                                  30'd    104    : data = 32'h    D45F8F93    ;    //    addi x31 x31 -699      ====        li x31, 0x1ad0bd45
                                                  30'd    105    : data = 32'h    800007B7    ;    //    lui x15 524288      ====        main: li a5, 0x80000000 #start riscv_int_numeric_corner_stream_10
                                                  30'd    106    : data = 32'h    00078793    ;    //    addi x15 x15 0      ====        main: li a5, 0x80000000 #start riscv_int_numeric_corner_stream_10
                                                  30'd    107    : data = 32'h    5A10D937    ;    //    lui x18 368909      ====        li s2, 0x5a10d661
                                                  30'd    108    : data = 32'h    66190913    ;    //    addi x18 x18 1633      ====        li s2, 0x5a10d661
                                                  30'd    109    : data = 32'h    FFF00413    ;    //    addi x8 x0 -1      ====        li s0, 0xffffffff
                                                  30'd    110    : data = 32'h    00000E93    ;    //    addi x29 x0 0      ====        li t4, 0x0
                                                  30'd    111    : data = 32'h    FFF00893    ;    //    addi x17 x0 -1      ====        li a7, 0xffffffff
                                                  30'd    112    : data = 32'h    35049CB7    ;    //    lui x25 217161      ====        li s9, 0x35049129
                                                  30'd    113    : data = 32'h    129C8C93    ;    //    addi x25 x25 297      ====        li s9, 0x35049129
                                                  30'd    114    : data = 32'h    FFF00393    ;    //    addi x7 x0 -1      ====        li t2, 0xffffffff
                                                  30'd    115    : data = 32'h    410546B7    ;    //    lui x13 266324      ====        li a3, 0x41053ec0
                                                  30'd    116    : data = 32'h    EC068693    ;    //    addi x13 x13 -320      ====        li a3, 0x41053ec0
                                                  30'd    117    : data = 32'h    D6124637    ;    //    lui x12 876836      ====        li a2, 0xd61247be
                                                  30'd    118    : data = 32'h    7BE60613    ;    //    addi x12 x12 1982      ====        li a2, 0xd61247be
                                                  30'd    119    : data = 32'h    BA354137    ;    //    lui x2 762708      ====        li sp, 0xba353e9c
                                                  30'd    120    : data = 32'h    E9C10113    ;    //    addi x2 x2 -356      ====        li sp, 0xba353e9c
                                                  30'd    121    : data = 32'h    01D78933    ;    //    add x18 x15 x29      ====        add s2, a5, t4
                                                  30'd    122    : data = 32'h    00C10133    ;    //    add x2 x2 x12      ====        add sp, sp, a2
                                                  30'd    123    : data = 32'h    007887B3    ;    //    add x15 x17 x7      ====        add a5, a7, t2
                                                  30'd    124    : data = 32'h    008908B3    ;    //    add x17 x18 x8      ====        add a7, s2, s0
                                                  30'd    125    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    126    : data = 32'h    412687B3    ;    //    sub x15 x13 x18      ====        sub a5, a3, s2
                                                  30'd    127    : data = 32'h    40288CB3    ;    //    sub x25 x17 x2      ====        sub s9, a7, sp
                                                  30'd    128    : data = 32'h    00F38EB3    ;    //    add x29 x7 x15      ====        add t4, t2, a5
                                                  30'd    129    : data = 32'h    8B8C8393    ;    //    addi x7 x25 -1864      ====        addi t2, s9, -1864
                                                  30'd    130    : data = 32'h    71FCDCB7    ;    //    lui x25 466893      ====        lui s9, 466893
                                                  30'd    131    : data = 32'h    61CE1E97    ;    //    auipc x29 400609      ====        auipc t4, 400609
                                                  30'd    132    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    133    : data = 32'h    4564DCB7    ;    //    lui x25 284237      ====        lui s9, 284237
                                                  30'd    134    : data = 32'h    01910EB3    ;    //    add x29 x2 x25      ====        add t4, sp, s9
                                                  30'd    135    : data = 32'h    00C90613    ;    //    addi x12 x18 12      ====        addi a2, s2, 12
                                                  30'd    136    : data = 32'h    92C4D117    ;    //    auipc x2 601165      ====        auipc sp, 601165
                                                  30'd    137    : data = 32'h    4AD40613    ;    //    addi x12 x8 1197      ====        addi a2, s0, 1197
                                                  30'd    138    : data = 32'h    40740CB3    ;    //    sub x25 x8 x7      ====        sub s9, s0, t2
                                                  30'd    139    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    140    : data = 32'h    A9E10917    ;    //    auipc x18 695824      ====        auipc s2, 695824
                                                  30'd    141    : data = 32'h    41938EB3    ;    //    sub x29 x7 x25      ====        sub t4, t2, s9
                                                  30'd    142    : data = 32'h    419608B3    ;    //    sub x17 x12 x25      ====        sub a7, a2, s9
                                                  30'd    143    : data = 32'h    BE888913    ;    //    addi x18 x17 -1048      ====        addi s2, a7, -1048
                                                  30'd    144    : data = 32'h    328D17B7    ;    //    lui x15 207057      ====        lui a5, 207057
                                                  30'd    145    : data = 32'h    7DD90113    ;    //    addi x2 x18 2013      ====        addi sp, s2, 2013
                                                  30'd    146    : data = 32'h    40C90633    ;    //    sub x12 x18 x12      ====        sub a2, s2, a2
                                                  30'd    147    : data = 32'h    8BF78893    ;    //    addi x17 x15 -1857      ====        addi a7, a5, -1857
                                                  30'd    148    : data = 32'h    41288EB3    ;    //    sub x29 x17 x18      ====        sub t4, a7, s2
                                                  30'd    149    : data = 32'h    0F8577B7    ;    //    lui x15 63575      ====        lui a5, 63575
                                                  30'd    150    : data = 32'h    407E87B3    ;    //    sub x15 x29 x7      ====        sub a5, t4, t2
                                               //   30'd    151    : data = 32'h    48C0B0EF    ;    //    jal  4x16220      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_10
                                                  30'd    152    : data = 32'h    800007B7    ;    //    lui x15 524288      ====        li a5, 0x80000000 #start riscv_int_numeric_corner_stream_22
                                                  30'd    153    : data = 32'h    00078793    ;    //    addi x15 x15 0      ====        li a5, 0x80000000 #start riscv_int_numeric_corner_stream_22
                                                  30'd    154    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff
                                                  30'd    155    : data = 32'h    FFF00293    ;    //    addi x5 x0 -1      ====        li t0, 0xffffffff
                                                  30'd    156    : data = 32'h    80000DB7    ;    //    lui x27 524288      ====        li s11, 0x80000000
                                                  30'd    157    : data = 32'h    000D8D93    ;    //    addi x27 x27 0      ====        li s11, 0x80000000
                                                  30'd    158    : data = 32'h    157C1A37    ;    //    lui x20 88001      ====        li s4, 0x157c126d
                                                  30'd    159    : data = 32'h    26DA0A13    ;    //    addi x20 x20 621      ====        li s4, 0x157c126d
                                                  30'd    160    : data = 32'h    80000D37    ;    //    lui x26 524288      ====        li s10, 0x80000000
                                                  30'd    161    : data = 32'h    000D0D13    ;    //    addi x26 x26 0      ====        li s10, 0x80000000
                                                  30'd    162    : data = 32'h    00000C13    ;    //    addi x24 x0 0      ====        li s8, 0x0
                                                  30'd    163    : data = 32'h    80000AB7    ;    //    lui x21 524288      ====        li s5, 0x80000000
                                                  30'd    164    : data = 32'h    000A8A93    ;    //    addi x21 x21 0      ====        li s5, 0x80000000
                                                  30'd    165    : data = 32'h    800006B7    ;    //    lui x13 524288      ====        li a3, 0x80000000
                                                  30'd    166    : data = 32'h    00068693    ;    //    addi x13 x13 0      ====        li a3, 0x80000000
                                                  30'd    167    : data = 32'h    00000193    ;    //    addi x3 x0 0      ====        li gp, 0x0
                                                  30'd    168    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    169    : data = 32'h    C2BF6D37    ;    //    lui x26 797686      ====        lui s10, 797686
                                                  30'd    170    : data = 32'h    403D06B3    ;    //    sub x13 x26 x3      ====        sub a3, s10, gp
                                                  30'd    171    : data = 32'h    1BBD0C13    ;    //    addi x24 x26 443      ====        addi s8, s10, 443
                                                  30'd    172    : data = 32'h    EF818797    ;    //    auipc x15 981016      ====        auipc a5, 981016
                                                  30'd    173    : data = 32'h    0DD28693    ;    //    addi x13 x5 221      ====        addi a3, t0, 221
                                                  30'd    174    : data = 32'h    00DD86B3    ;    //    add x13 x27 x13      ====        add a3, s11, a3
                                                  30'd    175    : data = 32'h    722D8A13    ;    //    addi x20 x27 1826      ====        addi s4, s11, 1826
                                                  30'd    176    : data = 32'h    9B00C797    ;    //    auipc x15 634892      ====        auipc a5, 634892
                                                  30'd    177    : data = 32'h    01878D33    ;    //    add x26 x15 x24      ====        add s10, a5, s8
                                                  30'd    178    : data = 32'h    CD9C0C13    ;    //    addi x24 x24 -807      ====        addi s8, s8, -807
                                                  30'd    179    : data = 32'h    9FD5B797    ;    //    auipc x15 654683      ====        auipc a5, 654683
                                                  30'd    180    : data = 32'h    5BBFC797    ;    //    auipc x15 375804      ====        auipc a5, 375804
                                                  30'd    181    : data = 32'h    F39D8D93    ;    //    addi x27 x27 -199      ====        addi s11, s11, -199
                                                  30'd    182    : data = 32'h    D24B5DB7    ;    //    lui x27 861365      ====        lui s11, 861365
                                                  30'd    183    : data = 32'h    C46A0D93    ;    //    addi x27 x20 -954      ====        addi s11, s4, -954
                                                  30'd    184    : data = 32'h    D2261AB7    ;    //    lui x21 860769      ====        lui s5, 860769
                                                  30'd    185    : data = 32'h    5C708C13    ;    //    addi x24 x1 1479      ====        addi s8, ra, 1479
                                                  30'd    186    : data = 32'h    CBB5F197    ;    //    auipc x3 834399      ====        auipc gp, 834399
                                                  30'd    187    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                              //    30'd    188    : data = 32'h    3F80B0EF    ;    //    jal x1 46072      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_22
                                                  30'd    189    : data = 32'h    2536AC37    ;    //    lui x24 152426      ====        li s8, 0x25369e12 #start riscv_int_numeric_corner_stream_4
                                                  30'd    190    : data = 32'h    E12C0C13    ;    //    addi x24 x24 -494      ====        li s8, 0x25369e12 #start riscv_int_numeric_corner_stream_4
                                                  30'd    191    : data = 32'h    65C67EB7    ;    //    lui x29 416871      ====        li t4, 0x65c66cfd
                                                  30'd    192    : data = 32'h    CFDE8E93    ;    //    addi x29 x29 -771      ====        li t4, 0x65c66cfd
                                                  30'd    193    : data = 32'h    00000E13    ;    //    addi x28 x0 0      ====        li t3, 0x0
                                                  30'd    194    : data = 32'h    FFF00993    ;    //    addi x19 x0 -1      ====        li s3, 0xffffffff
                                                  30'd    195    : data = 32'h    19059137    ;    //    lui x2 102489      ====        li sp, 0x190590fd
                                                  30'd    196    : data = 32'h    0FD10113    ;    //    addi x2 x2 253      ====        li sp, 0x190590fd
                                                  30'd    197    : data = 32'h    FFF00D13    ;    //    addi x26 x0 -1      ====        li s10, 0xffffffff
                                                  30'd    198    : data = 32'h    00000193    ;    //    addi x3 x0 0      ====        li gp, 0x0
                                                  30'd    199    : data = 32'h    F5E1A437    ;    //    lui x8 1007130      ====        li s0, 0xf5e1a1d6
                                                  30'd    200    : data = 32'h    1D640413    ;    //    addi x8 x8 470      ====        li s0, 0xf5e1a1d6
                                                  30'd    201    : data = 32'h    FFF00913    ;    //    addi x18 x0 -1      ====        li s2, 0xffffffff
                                                  30'd    202    : data = 32'h    0155C4B7    ;    //    lui x9 5468      ====        li s1, 0x155bc11
                                                  30'd    203    : data = 32'h    C1148493    ;    //    addi x9 x9 -1007      ====        li s1, 0x155bc11
                                                  30'd    204    : data = 32'h    408C0C33    ;    //    sub x24 x24 x8      ====        sub s8, s8, s0
                                                  30'd    205    : data = 32'h    3A540193    ;    //    addi x3 x8 933      ====        addi gp, s0, 933
                                                  30'd    206    : data = 32'h    E1E6D9B7    ;    //    lui x19 925293      ====        lui s3, 925293
                                                  30'd    207    : data = 32'h    B78D0193    ;    //    addi x3 x26 -1160      ====        addi gp, s10, -1160
                                                  30'd    208    : data = 32'h    009E8EB3    ;    //    add x29 x29 x9      ====        add t4, t4, s1
                                                  30'd    209    : data = 32'h    88B07137    ;    //    lui x2 559879      ====        lui sp, 559879
                                                  30'd    210    : data = 32'h    009E8933    ;    //    add x18 x29 x9      ====        add s2, t4, s1
                                                  30'd    211    : data = 32'h    41390433    ;    //    sub x8 x18 x19      ====        sub s0, s2, s3
                                                  30'd    212    : data = 32'h    F8CBD117    ;    //    auipc x2 1019069      ====        auipc sp, 1019069
                                                  30'd    213    : data = 32'h    41C18D33    ;    //    sub x26 x3 x28      ====        sub s10, gp, t3
                                                  30'd    214    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    215    : data = 32'h    00390133    ;    //    add x2 x18 x3      ====        add sp, s2, gp
                                                  30'd    216    : data = 32'h    FD018993    ;    //    addi x19 x3 -48      ====        addi s3, gp, -48
                                                  30'd    217    : data = 32'h    40840EB3    ;    //    sub x29 x8 x8      ====        sub t4, s0, s0
                                                  30'd    218    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    219    : data = 32'h    002E0E33    ;    //    add x28 x28 x2      ====        add t3, t3, sp
                                                  30'd    220    : data = 32'h    BD3D0D13    ;    //    addi x26 x26 -1069      ====        addi s10, s10, -1069
                                                  30'd    221    : data = 32'h    00840EB3    ;    //    add x29 x8 x8      ====        add t4, s0, s0
                                                  30'd    222    : data = 32'h    AB3E9C17    ;    //    auipc x24 701417      ====        auipc s8, 701417
                                                  30'd    223    : data = 32'h    37E51137    ;    //    lui x2 228945      ====        lui sp, 228945
                                                  30'd    224    : data = 32'h    A21AD937    ;    //    lui x18 663981      ====        lui s2, 663981
                                                  30'd    225    : data = 32'h    9DA24E17    ;    //    auipc x28 645668      ====        auipc t3, 645668
                                                  30'd    226    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    227    : data = 32'h    C99D7497    ;    //    auipc x9 825815      ====        auipc s1, 825815
                                                  30'd    228    : data = 32'h    1F740993    ;    //    addi x19 x8 503      ====        addi s3, s0, 503
                                                  30'd    229    : data = 32'h    91AB7137    ;    //    lui x2 596663      ====        lui sp, 596663
                                                  30'd    230    : data = 32'h    BCDC09B7    ;    //    lui x19 773568      ====        lui s3, 773568
                                                  30'd    231    : data = 32'h    95A98E13    ;    //    addi x28 x19 -1702      ====        addi t3, s3, -1702
                                                //  30'd    232    : data = 32'h    3480B0EF    ;    //    jal x1 45896      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_4
                                                  30'd    233    : data = 32'h    57B5DA37    ;    //    lui x20 359261      ====        li s4, 0x57b5c8c8 #start riscv_int_numeric_corner_stream_21
                                                  30'd    234    : data = 32'h    8C8A0A13    ;    //    addi x20 x20 -1848      ====        li s4, 0x57b5c8c8 #start riscv_int_numeric_corner_stream_21
                                                  30'd    235    : data = 32'h    800006B7    ;    //    lui x13 524288      ====        li a3, 0x80000000
                                                  30'd    236    : data = 32'h    00068693    ;    //    addi x13 x13 0      ====        li a3, 0x80000000
                                                  30'd    237    : data = 32'h    49E709B7    ;    //    lui x19 302704      ====        li s3, 0x49e6fb3e
                                                  30'd    238    : data = 32'h    B3E98993    ;    //    addi x19 x19 -1218      ====        li s3, 0x49e6fb3e
                                                  30'd    239    : data = 32'h    800001B7    ;    //    lui x3 524288      ====        li gp, 0x80000000
                                                  30'd    240    : data = 32'h    00018193    ;    //    addi x3 x3 0      ====        li gp, 0x80000000
                                                  30'd    241    : data = 32'h    FB4A5637    ;    //    lui x12 1029285      ====        li a2, 0xfb4a53f9
                                                  30'd    242    : data = 32'h    3F960613    ;    //    addi x12 x12 1017      ====        li a2, 0xfb4a53f9
                                                  30'd    243    : data = 32'h    80000CB7    ;    //    lui x25 524288      ====        li s9, 0x80000000
                                                  30'd    244    : data = 32'h    000C8C93    ;    //    addi x25 x25 0      ====        li s9, 0x80000000
                                                  30'd    245    : data = 32'h    FFF00A93    ;    //    addi x21 x0 -1      ====        li s5, 0xffffffff
                                                  30'd    246    : data = 32'h    FFF00F93    ;    //    addi x31 x0 -1      ====        li t6, 0xffffffff
                                                  30'd    247    : data = 32'h    80000E37    ;    //    lui x28 524288      ====        li t3, 0x80000000
                                                  30'd    248    : data = 32'h    000E0E13    ;    //    addi x28 x28 0      ====        li t3, 0x80000000
                                                  30'd    249    : data = 32'h    FFF00913    ;    //    addi x18 x0 -1      ====        li s2, 0xffffffff
                                                  30'd    250    : data = 32'h    419F8CB3    ;    //    sub x25 x31 x25      ====        sub s9, t6, s9
                                                  30'd    251    : data = 32'h    40DE01B3    ;    //    sub x3 x28 x13      ====        sub gp, t3, a3
                                                  30'd    252    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    253    : data = 32'h    00318CB3    ;    //    add x25 x3 x3      ====        add s9, gp, gp
                                                  30'd    254    : data = 32'h    A29B6697    ;    //    auipc x13 666038      ====        auipc a3, 666038
                                                  30'd    255    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    256    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    257    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    258    : data = 32'h    0279FC97    ;    //    auipc x25 10143      ====        auipc s9, 10143
                                                  30'd    259    : data = 32'h    59B12A97    ;    //    auipc x21 367378      ====        auipc s5, 367378
                                                  30'd    260    : data = 32'h    98494E37    ;    //    lui x28 623764      ====        lui t3, 623764
                                                  30'd    261    : data = 32'h    01F68933    ;    //    add x18 x13 x31      ====        add s2, a3, t6
                                                  30'd    262    : data = 32'h    415A8CB3    ;    //    sub x25 x21 x21      ====        sub s9, s5, s5
                                                  30'd    263    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    264    : data = 32'h    015981B3    ;    //    add x3 x19 x21      ====        add gp, s3, s5
                                                  30'd    265    : data = 32'h    40390A33    ;    //    sub x20 x18 x3      ====        sub s4, s2, gp
                                                  30'd    266    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    267    : data = 32'h    D1018693    ;    //    addi x13 x3 -752      ====        addi a3, gp, -752
                                                  30'd    268    : data = 32'h    C4990A93    ;    //    addi x21 x18 -951      ====        addi s5, s2, -951
                                                  30'd    269    : data = 32'h    212FF617    ;    //    auipc x12 135935      ====        auipc a2, 135935
                                                  30'd    270    : data = 32'h    A154B937    ;    //    lui x18 660811      ====        lui s2, 660811
                                               //   30'd    271    : data = 32'h    2AC0B0EF    ;    //    jal x1 45740      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_21
                                                  30'd    272    : data = 32'h    80000137    ;    //    lui x2 524288      ====        li sp, 0x80000000 #start riscv_int_numeric_corner_stream_29
                                                  30'd    273    : data = 32'h    00010113    ;    //    addi x2 x2 0      ====        li sp, 0x80000000 #start riscv_int_numeric_corner_stream_29
                                                  30'd    274    : data = 32'h    7BD0BBB7    ;    //    lui x23 507147      ====        li s7, 0x7bd0acfa
                                                  30'd    275    : data = 32'h    CFAB8B93    ;    //    addi x23 x23 -774      ====        li s7, 0x7bd0acfa
                                                  30'd    276    : data = 32'h    AF8E7CB7    ;    //    lui x25 719079      ====        li s9, 0xaf8e6f96
                                                  30'd    277    : data = 32'h    F96C8C93    ;    //    addi x25 x25 -106      ====        li s9, 0xaf8e6f96
                                                  30'd    278    : data = 32'h    FFF00593    ;    //    addi x11 x0 -1      ====        li a1, 0xffffffff
                                                  30'd    279    : data = 32'h    519FC4B7    ;    //    lui x9 334332      ====        li s1, 0x519fc133
                                                  30'd    280    : data = 32'h    13348493    ;    //    addi x9 x9 307      ====        li s1, 0x519fc133
                                                  30'd    281    : data = 32'h    80000837    ;    //    lui x16 524288      ====        li a6, 0x80000000
                                                  30'd    282    : data = 32'h    00080813    ;    //    addi x16 x16 0      ====        li a6, 0x80000000
                                                  30'd    283    : data = 32'h    F30058B7    ;    //    lui x17 995333      ====        li a7, 0xf300533f
                                                  30'd    284    : data = 32'h    33F88893    ;    //    addi x17 x17 831      ====        li a7, 0xf300533f
                                                  30'd    285    : data = 32'h    00000B13    ;    //    addi x22 x0 0      ====        li s6, 0x0
                                                  30'd    286    : data = 32'h    FFF00293    ;    //    addi x5 x0 -1      ====        li t0, 0xffffffff
                                                  30'd    287    : data = 32'h    FFF00A93    ;    //    addi x21 x0 -1      ====        li s5, 0xffffffff
                                                  30'd    288    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    289    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    290    : data = 32'h    DD080813    ;    //    addi x16 x16 -560      ====        addi a6, a6, -560
                                                  30'd    291    : data = 32'h    FE8574B7    ;    //    lui x9 1042519      ====        lui s1, 1042519
                                                  30'd    292    : data = 32'h    41780B33    ;    //    sub x22 x16 x23      ====        sub s6, a6, s7
                                                  30'd    293    : data = 32'h    010B02B3    ;    //    add x5 x22 x16      ====        add t0, s6, a6
                                                  30'd    294    : data = 32'h    40928133    ;    //    sub x2 x5 x9      ====        sub sp, t0, s1
                                                  30'd    295    : data = 32'h    B1F3FC97    ;    //    auipc x25 728895      ====        auipc s9, 728895
                                                  30'd    296    : data = 32'h    70D472B7    ;    //    lui x5 462151      ====        lui t0, 462151
                                                  30'd    297    : data = 32'h    AA428B93    ;    //    addi x23 x5 -1372      ====        addi s7, t0, -1372
                                                  30'd    298    : data = 32'h    CE258B93    ;    //    addi x23 x11 -798      ====        addi s7, a1, -798
                                                  30'd    299    : data = 32'h    B993D297    ;    //    auipc x5 760125      ====        auipc t0, 760125
                                                  30'd    300    : data = 32'h    409B02B3    ;    //    sub x5 x22 x9      ====        sub t0, s6, s1
                                                  30'd    301    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    302    : data = 32'h    11A58593    ;    //    addi x11 x11 282      ====        addi a1, a1, 282
                                                  30'd    303    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    304    : data = 32'h    010B0133    ;    //    add x2 x22 x16      ====        add sp, s6, a6
                                                  30'd    305    : data = 32'h    BA5A8813    ;    //    addi x16 x21 -1115      ====        addi a6, s5, -1115
                                                  30'd    306    : data = 32'h    40258133    ;    //    sub x2 x11 x2      ====        sub sp, a1, sp
                                                  30'd    307    : data = 32'h    01980BB3    ;    //    add x23 x16 x25      ====        add s7, a6, s9
                                                  30'd    308    : data = 32'h    40B805B3    ;    //    sub x11 x16 x11      ====        sub a1, a6, a1
                                                  30'd    309    : data = 32'h    CD242297    ;    //    auipc x5 840258      ====        auipc t0, 840258
                                               //   30'd    310    : data = 32'h    2100B0EF    ;    //    jal x1 45584      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_29
                                                  30'd    311    : data = 32'h    F84CB937    ;    //    lui x18 1017035      ====        li s2, 0xf84cb455 #start riscv_int_numeric_corner_stream_37
                                                  30'd    312    : data = 32'h    45590913    ;    //    addi x18 x18 1109      ====        li s2, 0xf84cb455 #start riscv_int_numeric_corner_stream_37
                                                  30'd    313    : data = 32'h    00000B93    ;    //    addi x23 x0 0      ====        li s7, 0x0
                                                  30'd    314    : data = 32'h    12EFF2B7    ;    //    lui x5 77567      ====        li t0, 0x12efedab
                                                  30'd    315    : data = 32'h    DAB28293    ;    //    addi x5 x5 -597      ====        li t0, 0x12efedab
                                                  30'd    316    : data = 32'h    0D01A4B7    ;    //    lui x9 53274      ====        li s1, 0xd01a71b
                                                  30'd    317    : data = 32'h    71B48493    ;    //    addi x9 x9 1819      ====        li s1, 0xd01a71b
                                                  30'd    318    : data = 32'h    BC994D37    ;    //    lui x26 772500      ====        li s10, 0xbc993d4f
                                                  30'd    319    : data = 32'h    D4FD0D13    ;    //    addi x26 x26 -689      ====        li s10, 0xbc993d4f
                                                  30'd    320    : data = 32'h    00000713    ;    //    addi x14 x0 0      ====        li a4, 0x0
                                                  30'd    321    : data = 32'h    FFF00413    ;    //    addi x8 x0 -1      ====        li s0, 0xffffffff
                                                  30'd    322    : data = 32'h    80000A37    ;    //    lui x20 524288      ====        li s4, 0x80000000
                                                  30'd    323    : data = 32'h    000A0A13    ;    //    addi x20 x20 0      ====        li s4, 0x80000000
                                                  30'd    324    : data = 32'h    FFF00893    ;    //    addi x17 x0 -1      ====        li a7, 0xffffffff
                                                  30'd    325    : data = 32'h    5D1D73B7    ;    //    lui x7 381399      ====        li t2, 0x5d1d74a4
                                                  30'd    326    : data = 32'h    4A438393    ;    //    addi x7 x7 1188      ====        li t2, 0x5d1d74a4
                                                  30'd    327    : data = 32'h    5B237B97    ;    //    auipc x23 373303      ====        auipc s7, 373303
                                                  30'd    328    : data = 32'h    012288B3    ;    //    add x17 x5 x18      ====        add a7, t0, s2
                                                  30'd    329    : data = 32'h    40E40A33    ;    //    sub x20 x8 x14      ====        sub s4, s0, a4
                                                  30'd    330    : data = 32'h    01AD03B3    ;    //    add x7 x26 x26      ====        add t2, s10, s10
                                                  30'd    331    : data = 32'h    CC048293    ;    //    addi x5 x9 -832      ====        addi t0, s1, -832
                                                  30'd    332    : data = 32'h    6B6A2737    ;    //    lui x14 439970      ====        lui a4, 439970
                                                  30'd    333    : data = 32'h    BED70B93    ;    //    addi x23 x14 -1043      ====        addi s7, a4, -1043
                                                  30'd    334    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    335    : data = 32'h    7AF20717    ;    //    auipc x14 503584      ====        auipc a4, 503584
                                                  30'd    336    : data = 32'h    007404B3    ;    //    add x9 x8 x7      ====        add s1, s0, t2
                                                  30'd    337    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    338    : data = 32'h    0E8A0B93    ;    //    addi x23 x20 232      ====        addi s7, s4, 232
                                                  30'd    339    : data = 32'h    6AC86397    ;    //    auipc x7 437382      ====        auipc t2, 437382
                                                  30'd    340    : data = 32'h    412883B3    ;    //    sub x7 x17 x18      ====        sub t2, a7, s2
                                                  30'd    341    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    342    : data = 32'h    017404B3    ;    //    add x9 x8 x23      ====        add s1, s0, s7
                                                  30'd    343    : data = 32'h    7400C297    ;    //    auipc x5 475148      ====        auipc t0, 475148
                                                  30'd    344    : data = 32'h    40928433    ;    //    sub x8 x5 x9      ====        sub s0, t0, s1
                                                  30'd    345    : data = 32'h    4C387737    ;    //    lui x14 312199      ====        lui a4, 312199
                                                  30'd    346    : data = 32'h    786984B7    ;    //    lui x9 493208      ====        lui s1, 493208
                                                  30'd    347    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    348    : data = 32'h    0096B297    ;    //    auipc x5 2411      ====        auipc t0, 2411
                                                  30'd    349    : data = 32'h    A2712417    ;    //    auipc x8 665362      ====        auipc s0, 665362
                                               //   30'd    350    : data = 32'h    1700B0EF    ;    //    jal x1 45424      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_37
                                                  30'd    351    : data = 32'h    45FA2337    ;    //    lui x6 286626      ====        li t1, 0x45fa2248 #start riscv_int_numeric_corner_stream_24
                                                  30'd    352    : data = 32'h    24830313    ;    //    addi x6 x6 584      ====        li t1, 0x45fa2248 #start riscv_int_numeric_corner_stream_24
                                                  30'd    353    : data = 32'h    80000AB7    ;    //    lui x21 524288      ====        li s5, 0x80000000
                                                  30'd    354    : data = 32'h    000A8A93    ;    //    addi x21 x21 0      ====        li s5, 0x80000000
                                                  30'd    355    : data = 32'h    00000393    ;    //    addi x7 x0 0      ====        li t2, 0x0
                                                  30'd    356    : data = 32'h    220C0937    ;    //    lui x18 139456      ====        li s2, 0x220bf84d
                                                  30'd    357    : data = 32'h    84D90913    ;    //    addi x18 x18 -1971      ====        li s2, 0x220bf84d
                                                  30'd    358    : data = 32'h    00000093    ;    //    addi x1 x0 0      ====        li ra, 0x0
                                                  30'd    359    : data = 32'h    FFF00113    ;    //    addi x2 x0 -1      ====        li sp, 0xffffffff
                                                  30'd    360    : data = 32'h    FFF00613    ;    //    addi x12 x0 -1      ====        li a2, 0xffffffff
                                                  30'd    361    : data = 32'h    E78C6EB7    ;    //    lui x29 948422      ====        li t4, 0xe78c6534
                                                  30'd    362    : data = 32'h    534E8E93    ;    //    addi x29 x29 1332      ====        li t4, 0xe78c6534
                                                  30'd    363    : data = 32'h    FE598B37    ;    //    lui x22 1041816      ====        li s6, 0xfe597c60
                                                  30'd    364    : data = 32'h    C60B0B13    ;    //    addi x22 x22 -928      ====        li s6, 0xfe597c60
                                                  30'd    365    : data = 32'h    FFF00193    ;    //    addi x3 x0 -1      ====        li gp, 0xffffffff
                                                  30'd    366    : data = 32'h    74810093    ;    //    addi x1 x2 1864      ====        addi ra, sp, 1864
                                                  30'd    367    : data = 32'h    007101B3    ;    //    add x3 x2 x7      ====        add gp, sp, t2
                                                  30'd    368    : data = 32'h    C41F9637    ;    //    lui x12 803321      ====        lui a2, 803321
                                                  30'd    369    : data = 32'h    685B0E93    ;    //    addi x29 x22 1669      ====        addi t4, s6, 1669
                                                  30'd    370    : data = 32'h    01DB0633    ;    //    add x12 x22 x29      ====        add a2, s6, t4
                                                  30'd    371    : data = 32'h    3E81E617    ;    //    auipc x12 256030      ====        auipc a2, 256030
                                                  30'd    372    : data = 32'h    006100B3    ;    //    add x1 x2 x6      ====        add ra, sp, t1
                                                  30'd    373    : data = 32'h    00760633    ;    //    add x12 x12 x7      ====        add a2, a2, t2
                                                  30'd    374    : data = 32'h    2D290913    ;    //    addi x18 x18 722      ====        addi s2, s2, 722
                                                  30'd    375    : data = 32'h    00160933    ;    //    add x18 x12 x1      ====        add s2, a2, ra
                                                  30'd    376    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    377    : data = 32'h    8A03EAB7    ;    //    lui x21 565310      ====        lui s5, 565310
                                                  30'd    378    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    379    : data = 32'h    2B4B0193    ;    //    addi x3 x22 692      ====        addi gp, s6, 692
                                                  30'd    380    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    381    : data = 32'h    002A8B33    ;    //    add x22 x21 x2      ====        add s6, s5, sp
                                                  30'd    382    : data = 32'h    01530633    ;    //    add x12 x6 x21      ====        add a2, t1, s5
                                                  30'd    383    : data = 32'h    41627E97    ;    //    auipc x29 267815      ====        auipc t4, 267815
                                                  30'd    384    : data = 32'h    B1EC8637    ;    //    lui x12 728776      ====        lui a2, 728776
                                                  30'd    385    : data = 32'h    01260933    ;    //    add x18 x12 x18      ====        add s2, a2, s2
                                                  30'd    386    : data = 32'h    1C6E8113    ;    //    addi x2 x29 454      ====        addi sp, t4, 454
                                                  30'd    387    : data = 32'h    1DC75B37    ;    //    lui x22 121973      ====        lui s6, 121973
                                                  30'd    388    : data = 32'h    36DD2937    ;    //    lui x18 224722      ====        lui s2, 224722
                                                  30'd    389    : data = 32'h    78156317    ;    //    auipc x6 491862      ====        auipc t1, 491862
                                                  30'd    390    : data = 32'h    41D30AB3    ;    //    sub x21 x6 x29      ====        sub s5, t1, t4
                                                  30'd    391    : data = 32'h    00338633    ;    //    add x12 x7 x3      ====        add a2, t2, gp
                                                  30'd    392    : data = 32'h    888B0093    ;    //    addi x1 x22 -1912      ====        addi ra, s6, -1912
                                                  30'd    393    : data = 32'h    40760B33    ;    //    sub x22 x12 x7      ====        sub s6, a2, t2
                                                //  30'd    394    : data = 32'h    0C00B0EF    ;    //    jal x1 45248      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_24
                                                  30'd    395    : data = 32'h    80000EB7    ;    //    lui x29 524288      ====        li t4, 0x80000000 #start riscv_int_numeric_corner_stream_27
                                                  30'd    396    : data = 32'h    000E8E93    ;    //    addi x29 x29 0      ====        li t4, 0x80000000 #start riscv_int_numeric_corner_stream_27
                                                  30'd    397    : data = 32'h    D3F4B4B7    ;    //    lui x9 868171      ====        li s1, 0xd3f4aa26
                                                  30'd    398    : data = 32'h    A2648493    ;    //    addi x9 x9 -1498      ====        li s1, 0xd3f4aa26
                                                  30'd    399    : data = 32'h    0B6F10B7    ;    //    lui x1 46833      ====        li ra, 0xb6f12e8
                                                  30'd    400    : data = 32'h    2E808093    ;    //    addi x1 x1 744      ====        li ra, 0xb6f12e8
                                                  30'd    401    : data = 32'h    F7A553B7    ;    //    lui x7 1014357      ====        li t2, 0xf7a555ad
                                                  30'd    402    : data = 32'h    5AD38393    ;    //    addi x7 x7 1453      ====        li t2, 0xf7a555ad
                                                  30'd    403    : data = 32'h    80000CB7    ;    //    lui x25 524288      ====        li s9, 0x80000000
                                                  30'd    404    : data = 32'h    000C8C93    ;    //    addi x25 x25 0      ====        li s9, 0x80000000
                                                  30'd    405    : data = 32'h    FFF00F93    ;    //    addi x31 x0 -1      ====        li t6, 0xffffffff
                                                  30'd    406    : data = 32'h    00000593    ;    //    addi x11 x0 0      ====        li a1, 0x0
                                                  30'd    407    : data = 32'h    FFF00293    ;    //    addi x5 x0 -1      ====        li t0, 0xffffffff
                                                  30'd    408    : data = 32'h    00000713    ;    //    addi x14 x0 0      ====        li a4, 0x0
                                                  30'd    409    : data = 32'h    E991B137    ;    //    lui x2 956699      ====        li sp, 0xe991a96c
                                                  30'd    410    : data = 32'h    96C10113    ;    //    addi x2 x2 -1684      ====        li sp, 0xe991a96c
                                                  30'd    411    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    412    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    413    : data = 32'h    40710FB3    ;    //    sub x31 x2 x7      ====        sub t6, sp, t2
                                                  30'd    414    : data = 32'h    B3D5B0B7    ;    //    lui x1 736603      ====        lui ra, 736603
                                                  30'd    415    : data = 32'h    409F8733    ;    //    sub x14 x31 x9      ====        sub a4, t6, s1
                                                  30'd    416    : data = 32'h    F0E38713    ;    //    addi x14 x7 -242      ====        addi a4, t2, -242
                                                  30'd    417    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    418    : data = 32'h    40B583B3    ;    //    sub x7 x11 x11      ====        sub t2, a1, a1
                                                  30'd    419    : data = 32'h    DB110493    ;    //    addi x9 x2 -591      ====        addi s1, sp, -591
                                                  30'd    420    : data = 32'h    56228C93    ;    //    addi x25 x5 1378      ====        addi s9, t0, 1378
                                                  30'd    421    : data = 32'h    D8CA5137    ;    //    lui x2 887973      ====        lui sp, 887973
                                                  30'd    422    : data = 32'h    FF80C397    ;    //    auipc x7 1046540      ====        auipc t2, 1046540
                                                  30'd    423    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    424    : data = 32'h    00E385B3    ;    //    add x11 x7 x14      ====        add a1, t2, a4
                                                  30'd    425    : data = 32'h    C0A44737    ;    //    lui x14 789060      ====        lui a4, 789060
                                                  30'd    426    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    427    : data = 32'h    6A0B2737    ;    //    lui x14 434354      ====        lui a4, 434354
                                                  30'd    428    : data = 32'h    278800B7    ;    //    lui x1 161920      ====        lui ra, 161920
                                                  30'd    429    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    430    : data = 32'h    D9C38C93    ;    //    addi x25 x7 -612      ====        addi s9, t2, -612
                                                  30'd    431    : data = 32'h    A9EE1EB7    ;    //    lui x29 696033      ====        lui t4, 696033
                                                  30'd    432    : data = 32'h    40E10133    ;    //    sub x2 x2 x14      ====        sub sp, sp, a4
                                                  30'd    433    : data = 32'h    F7571137    ;    //    lui x2 1013105      ====        lui sp, 1013105
                                                  30'd    434    : data = 32'h    2D138F93    ;    //    addi x31 x7 721      ====        addi t6, t2, 721
                                                  30'd    435    : data = 32'h    22D64597    ;    //    auipc x11 142692      ====        auipc a1, 142692
                                               //   30'd    436    : data = 32'h    0180B0EF    ;    //    jal x1 45080      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_27
                                                  30'd    437    : data = 32'h    FFF00393    ;    //    addi x7 x0 -1      ====        li t2, 0xffffffff #start riscv_int_numeric_corner_stream_39
                                                  30'd    438    : data = 32'h    38D299B7    ;    //    lui x19 232745      ====        li s3, 0x38d2979d
                                                  30'd    439    : data = 32'h    79D98993    ;    //    addi x19 x19 1949      ====        li s3, 0x38d2979d
                                                  30'd    440    : data = 32'h    00000A93    ;    //    addi x21 x0 0      ====        li s5, 0x0
                                                  30'd    441    : data = 32'h    00000593    ;    //    addi x11 x0 0      ====        li a1, 0x0
                                                  30'd    442    : data = 32'h    00000E13    ;    //    addi x28 x0 0      ====        li t3, 0x0
                                                  30'd    443    : data = 32'h    FFF00413    ;    //    addi x8 x0 -1      ====        li s0, 0xffffffff
                                                  30'd    444    : data = 32'h    80000137    ;    //    lui x2 524288      ====        li sp, 0x80000000
                                                  30'd    445    : data = 32'h    00010113    ;    //    addi x2 x2 0      ====        li sp, 0x80000000
                                                  30'd    446    : data = 32'h    00000893    ;    //    addi x17 x0 0      ====        li a7, 0x0
                                                  30'd    447    : data = 32'h    00000313    ;    //    addi x6 x0 0      ====        li t1, 0x0
                                                  30'd    448    : data = 32'h    FFF00293    ;    //    addi x5 x0 -1      ====        li t0, 0xffffffff
                                                  30'd    449    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    450    : data = 32'h    7510B9B7    ;    //    lui x19 479499      ====        lui s3, 479499
                                                  30'd    451    : data = 32'h    899EB997    ;    //    auipc x19 563691      ====        auipc s3, 563691
                                                  30'd    452    : data = 32'h    40B30433    ;    //    sub x8 x6 x11      ====        sub s0, t1, a1
                                                  30'd    453    : data = 32'h    CAB91997    ;    //    auipc x19 830353      ====        auipc s3, 830353
                                                  30'd    454    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    455    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    456    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    457    : data = 32'h    52AA1437    ;    //    lui x8 338593      ====        lui s0, 338593
                                                  30'd    458    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    459    : data = 32'h    FFCA8E13    ;    //    addi x28 x21 -4      ====        addi t3, s5, -4
                                                  30'd    460    : data = 32'h    013302B3    ;    //    add x5 x6 x19      ====        add t0, t1, s3
                                                  30'd    461    : data = 32'h    EC0E8297    ;    //    auipc x5 966888      ====        auipc t0, 966888
                                                  30'd    462    : data = 32'h    05784997    ;    //    auipc x19 22404      ====        auipc s3, 22404
                                                  30'd    463    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    464    : data = 32'h    005583B3    ;    //    add x7 x11 x5      ====        add t2, a1, t0
                                                  30'd    465    : data = 32'h    40630333    ;    //    sub x6 x6 x6      ====        sub t1, t1, t1
                                                  30'd    466    : data = 32'h    406288B3    ;    //    sub x17 x5 x6      ====        sub a7, t0, t1
                                                  30'd    467    : data = 32'h    4751B2B7    ;    //    lui x5 292123      ====        lui t0, 292123
                                                  30'd    468    : data = 32'h    AF030593    ;    //    addi x11 x6 -1296      ====        addi a1, t1, -1296
                                                  30'd    469    : data = 32'h    406E0433    ;    //    sub x8 x28 x6      ====        sub s0, t3, t1
                                                  30'd    470    : data = 32'h    413303B3    ;    //    sub x7 x6 x19      ====        sub t2, t1, s3
                                                  30'd    471    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    472    : data = 32'h    AF358593    ;    //    addi x11 x11 -1293      ====        addi a1, a1, -1293
                                                  30'd    473    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    474    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    475    : data = 32'h    007582B3    ;    //    add x5 x11 x7      ====        add t0, a1, t2
                                                  30'd    476    : data = 32'h    DC640413    ;    //    addi x8 x8 -570      ====        addi s0, s0, -570
                                               //   30'd    477    : data = 32'h    7750A0EF    ;    //    jal x1 44916      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_39
                                                  30'd    478    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff #start riscv_int_numeric_corner_stream_9
                                                  30'd    479    : data = 32'h    80000137    ;    //    lui x2 524288      ====        li sp, 0x80000000
                                                  30'd    480    : data = 32'h    00010113    ;    //    addi x2 x2 0      ====        li sp, 0x80000000
                                                  30'd    481    : data = 32'h    00000C13    ;    //    addi x24 x0 0      ====        li s8, 0x0
                                                  30'd    482    : data = 32'h    FFF00A93    ;    //    addi x21 x0 -1      ====        li s5, 0xffffffff
                                                  30'd    483    : data = 32'h    80000B37    ;    //    lui x22 524288      ====        li s6, 0x80000000
                                                  30'd    484    : data = 32'h    000B0B13    ;    //    addi x22 x22 0      ====        li s6, 0x80000000
                                                  30'd    485    : data = 32'h    FFF00C93    ;    //    addi x25 x0 -1      ====        li s9, 0xffffffff
                                                  30'd    486    : data = 32'h    00000393    ;    //    addi x7 x0 0      ====        li t2, 0x0
                                                  30'd    487    : data = 32'h    FFF00B93    ;    //    addi x23 x0 -1      ====        li s7, 0xffffffff
                                                  30'd    488    : data = 32'h    80000637    ;    //    lui x12 524288      ====        li a2, 0x80000000
                                                  30'd    489    : data = 32'h    00060613    ;    //    addi x12 x12 0      ====        li a2, 0x80000000
                                                  30'd    490    : data = 32'h    55B2D5B7    ;    //    lui x11 351021      ====        li a1, 0x55b2ccfe
                                                  30'd    491    : data = 32'h    CFE58593    ;    //    addi x11 x11 -770      ====        li a1, 0x55b2ccfe
                                                  30'd    492    : data = 32'h    47BA2637    ;    //    lui x12 293794      ====        lui a2, 293794
                                                  30'd    493    : data = 32'h    E3463BB7    ;    //    lui x23 930915      ====        lui s7, 930915
                                                  30'd    494    : data = 32'h    002B0CB3    ;    //    add x25 x22 x2      ====        add s9, s6, sp
                                                  30'd    495    : data = 32'h    DC4D25B7    ;    //    lui x11 902354      ====        lui a1, 902354
                                                  30'd    496    : data = 32'h    F8C27117    ;    //    auipc x2 1018919      ====        auipc sp, 1018919
                                                  30'd    497    : data = 32'h    017385B3    ;    //    add x11 x7 x23      ====        add a1, t2, s7
                                                  30'd    498    : data = 32'h    9DA10A93    ;    //    addi x21 x2 -1574      ====        addi s5, sp, -1574
                                                  30'd    499    : data = 32'h    01960CB3    ;    //    add x25 x12 x25      ====        add s9, a2, s9
                                                  30'd    500    : data = 32'h    F2B0B0B7    ;    //    lui x1 994059      ====        lui ra, 994059
                                                  30'd    501    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    502    : data = 32'h    6D7AACB7    ;    //    lui x25 448426      ====        lui s9, 448426
                                                  30'd    503    : data = 32'h    CF938A93    ;    //    addi x21 x7 -775      ====        addi s5, t2, -775
                                                  30'd    504    : data = 32'h    419C80B3    ;    //    sub x1 x25 x25      ====        sub ra, s9, s9
                                                  30'd    505    : data = 32'h    21712397    ;    //    auipc x7 136978      ====        auipc t2, 136978
                                                  30'd    506    : data = 32'h    40C38AB3    ;    //    sub x21 x7 x12      ====        sub s5, t2, a2
                                                  30'd    507    : data = 32'h    00CB0133    ;    //    add x2 x22 x12      ====        add sp, s6, a2
                                                  30'd    508    : data = 32'h    01958633    ;    //    add x12 x11 x25      ====        add a2, a1, s9
                                                  30'd    509    : data = 32'h    86308C13    ;    //    addi x24 x1 -1949      ====        addi s8, ra, -1949
                                                  30'd    510    : data = 32'h    872B0613    ;    //    addi x12 x22 -1934      ====        addi a2, s6, -1934
                                                  30'd    511    : data = 32'h    2BB635B7    ;    //    lui x11 179043      ====        lui a1, 179043
                                                  30'd    512    : data = 32'h    33D25B37    ;    //    lui x22 212261      ====        lui s6, 212261
                                                  30'd    513    : data = 32'h    CCDE9137    ;    //    lui x2 839145      ====        lui sp, 839145
                                                  30'd    514    : data = 32'h    00BB8633    ;    //    add x12 x23 x11      ====        add a2, s7, a1
                                                  30'd    515    : data = 32'h    01658B33    ;    //    add x22 x11 x22      ====        add s6, a1, s6
                                                  30'd    516    : data = 32'h    82E6BA97    ;    //    auipc x21 536171      ====        auipc s5, 536171
                                                  30'd    517    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    518    : data = 32'h    415C8633    ;    //    sub x12 x25 x21      ====        sub a2, s9, s5
                                                  30'd    519    : data = 32'h    8520CC97    ;    //    auipc x25 545292      ====        auipc s9, 545292
                                                  30'd    520    : data = 32'h    B782C5B7    ;    //    lui x11 751660      ====        lui a1, 751660
                                                //  30'd    521    : data = 32'h    6C50A0EF    ;    //    jal x1 44740      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_9
                                                  30'd    522    : data = 32'h    33525437    ;    //    lui x8 210213      ====        li s0, 0x335253fa #start riscv_int_numeric_corner_stream_26
                                                  30'd    523    : data = 32'h    3FA40413    ;    //    addi x8 x8 1018      ====        li s0, 0x335253fa #start riscv_int_numeric_corner_stream_26
                                                  30'd    524    : data = 32'h    FFF00713    ;    //    addi x14 x0 -1      ====        li a4, 0xffffffff
                                                  30'd    525    : data = 32'h    80000DB7    ;    //    lui x27 524288      ====        li s11, 0x80000000
                                                  30'd    526    : data = 32'h    000D8D93    ;    //    addi x27 x27 0      ====        li s11, 0x80000000
                                                  30'd    527    : data = 32'h    C88AF7B7    ;    //    lui x15 821423      ====        li a5, 0xc88af75b
                                                  30'd    528    : data = 32'h    75B78793    ;    //    addi x15 x15 1883      ====        li a5, 0xc88af75b
                                                  30'd    529    : data = 32'h    FFF00993    ;    //    addi x19 x0 -1      ====        li s3, 0xffffffff
                                                  30'd    530    : data = 32'h    800005B7    ;    //    lui x11 524288      ====        li a1, 0x80000000
                                                  30'd    531    : data = 32'h    00058593    ;    //    addi x11 x11 0      ====        li a1, 0x80000000
                                                  30'd    532    : data = 32'h    FFF00B93    ;    //    addi x23 x0 -1      ====        li s7, 0xffffffff
                                                  30'd    533    : data = 32'h    DDD15A37    ;    //    lui x20 908565      ====        li s4, 0xddd1523c
                                                  30'd    534    : data = 32'h    23CA0A13    ;    //    addi x20 x20 572      ====        li s4, 0xddd1523c
                                                  30'd    535    : data = 32'h    FFF00A93    ;    //    addi x21 x0 -1      ====        li s5, 0xffffffff
                                                  30'd    536    : data = 32'h    E8DF9D37    ;    //    lui x26 953849      ====        li s10, 0xe8df8e05
                                                  30'd    537    : data = 32'h    E05D0D13    ;    //    addi x26 x26 -507      ====        li s10, 0xe8df8e05
                                                  30'd    538    : data = 32'h    40BA0BB3    ;    //    sub x23 x20 x11      ====        sub s7, s4, a1
                                                  30'd    539    : data = 32'h    346B8593    ;    //    addi x11 x23 838      ====        addi a1, s7, 838
                                                  30'd    540    : data = 32'h    01AB8D33    ;    //    add x26 x23 x26      ====        add s10, s7, s10
                                                  30'd    541    : data = 32'h    103A8993    ;    //    addi x19 x21 259      ====        addi s3, s5, 259
                                                  30'd    542    : data = 32'h    A9718A17    ;    //    auipc x20 694040      ====        auipc s4, 694040
                                                  30'd    543    : data = 32'h    014A0BB3    ;    //    add x23 x20 x20      ====        add s7, s4, s4
                                                  30'd    544    : data = 32'h    40F78733    ;    //    sub x14 x15 x15      ====        sub a4, a5, a5
                                                  30'd    545    : data = 32'h    5F978D13    ;    //    addi x26 x15 1529      ====        addi s10, a5, 1529
                                                  30'd    546    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    547    : data = 32'h    CA6C4D97    ;    //    auipc x27 829124      ====        auipc s11, 829124
                                                  30'd    548    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    549    : data = 32'h    00EA0433    ;    //    add x8 x20 x14      ====        add s0, s4, a4
                                                  30'd    550    : data = 32'h    59DD5D37    ;    //    lui x26 368085      ====        lui s10, 368085
                                                  30'd    551    : data = 32'h    75A78713    ;    //    addi x14 x15 1882      ====        addi a4, a5, 1882
                                                  30'd    552    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    553    : data = 32'h    A981B5B7    ;    //    lui x11 694299      ====        lui a1, 694299
                                                  30'd    554    : data = 32'h    417B8A33    ;    //    sub x20 x23 x23      ====        sub s4, s7, s7
                                                  30'd    555    : data = 32'h    40840AB3    ;    //    sub x21 x8 x8      ====        sub s5, s0, s0
                                                  30'd    556    : data = 32'h    0C758713    ;    //    addi x14 x11 199      ====        addi a4, a1, 199
                                                  30'd    557    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    558    : data = 32'h    0D9D1417    ;    //    auipc x8 55761      ====        auipc s0, 55761
                                                  30'd    559    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    560    : data = 32'h    413D8DB3    ;    //    sub x27 x27 x19      ====        sub s11, s11, s3
                                                  30'd    561    : data = 32'h    01458433    ;    //    add x8 x11 x20      ====        add s0, a1, s4
                                                  30'd    562    : data = 32'h    F6B7DD17    ;    //    auipc x26 1010557      ====        auipc s10, 1010557
                                                  30'd    563    : data = 32'h    A0ADDD37    ;    //    lui x26 658141      ====        lui s10, 658141
                                                  30'd    564    : data = 32'h    40B98733    ;    //    sub x14 x19 x11      ====        sub a4, s3, a1
                                                  30'd    565    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    566    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    567    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                 // 30'd    568    : data = 32'h    6090A0EF    ;    //    jal x1 44552      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_26
                                                  30'd    569    : data = 32'h    00000113    ;    //    addi x2 x0 0      ====        li sp, 0x0 #start riscv_int_numeric_corner_stream_6
                                                  30'd    570    : data = 32'h    AE9BF4B7    ;    //    lui x9 715199      ====        li s1, 0xae9bf065
                                                  30'd    571    : data = 32'h    06548493    ;    //    addi x9 x9 101      ====        li s1, 0xae9bf065
                                                  30'd    572    : data = 32'h    446D16B7    ;    //    lui x13 280273      ====        li a3, 0x446d0933
                                                  30'd    573    : data = 32'h    93368693    ;    //    addi x13 x13 -1741      ====        li a3, 0x446d0933
                                                  30'd    574    : data = 32'h    00000C93    ;    //    addi x25 x0 0      ====        li s9, 0x0
                                                  30'd    575    : data = 32'h    00000193    ;    //    addi x3 x0 0      ====        li gp, 0x0
                                                  30'd    576    : data = 32'h    FFF00B13    ;    //    addi x22 x0 -1      ====        li s6, 0xffffffff
                                                  30'd    577    : data = 32'h    B4B72FB7    ;    //    lui x31 740210      ====        li t6, 0xb4b71a5b
                                                  30'd    578    : data = 32'h    A5BF8F93    ;    //    addi x31 x31 -1445      ====        li t6, 0xb4b71a5b
                                                  30'd    579    : data = 32'h    800000B7    ;    //    lui x1 524288      ====        li ra, 0x80000000
                                                  30'd    580    : data = 32'h    00008093    ;    //    addi x1 x1 0      ====        li ra, 0x80000000
                                                  30'd    581    : data = 32'h    80000937    ;    //    lui x18 524288      ====        li s2, 0x80000000
                                                  30'd    582    : data = 32'h    00090913    ;    //    addi x18 x18 0      ====        li s2, 0x80000000
                                                  30'd    583    : data = 32'h    98D19E37    ;    //    lui x28 625945      ====        li t3, 0x98d191a8
                                                  30'd    584    : data = 32'h    1A8E0E13    ;    //    addi x28 x28 424      ====        li t3, 0x98d191a8
                                                  30'd    585    : data = 32'h    001484B3    ;    //    add x9 x9 x1      ====        add s1, s1, ra
                                                  30'd    586    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    587    : data = 32'h    3EE58B17    ;    //    auipc x22 257624      ====        auipc s6, 257624
                                                  30'd    588    : data = 32'h    A3F0BB37    ;    //    lui x22 671499      ====        lui s6, 671499
                                                  30'd    589    : data = 32'h    87CA2F97    ;    //    auipc x31 556194      ====        auipc t6, 556194
                                                  30'd    590    : data = 32'h    419E0E33    ;    //    sub x28 x28 x25      ====        sub t3, t3, s9
                                                  30'd    591    : data = 32'h    C8963F97    ;    //    auipc x31 821603      ====        auipc t6, 821603
                                                  30'd    592    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    593    : data = 32'h    33EF8E13    ;    //    addi x28 x31 830      ====        addi t3, t6, 830
                                                  30'd    594    : data = 32'h    E6555E17    ;    //    auipc x28 943445      ====        auipc t3, 943445
                                                  30'd    595    : data = 32'h    9F8ECB17    ;    //    auipc x22 653548      ====        auipc s6, 653548
                                                  30'd    596    : data = 32'h    BFC71197    ;    //    auipc x3 785521      ====        auipc gp, 785521
                                                  30'd    597    : data = 32'h    001086B3    ;    //    add x13 x1 x1      ====        add a3, ra, ra
                                                  30'd    598    : data = 32'h    97F4DE37    ;    //    lui x28 622413      ====        lui t3, 622413
                                                  30'd    599    : data = 32'h    73E68937    ;    //    lui x18 474728      ====        lui s2, 474728
                                                 // 30'd    600    : data = 32'h    5890A0EF    ;    //    jal x1 44424      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_6
                                                  30'd    601    : data = 32'h    00000693    ;    //    addi x13 x0 0      ====        li a3, 0x0 #start riscv_int_numeric_corner_stream_20
                                                  30'd    602    : data = 32'h    00000193    ;    //    addi x3 x0 0      ====        li gp, 0x0
                                                  30'd    603    : data = 32'h    17826637    ;    //    lui x12 96294      ====        li a2, 0x17825de0
                                                  30'd    604    : data = 32'h    DE060613    ;    //    addi x12 x12 -544      ====        li a2, 0x17825de0
                                                  30'd    605    : data = 32'h    00000913    ;    //    addi x18 x0 0      ====        li s2, 0x0
                                                  30'd    606    : data = 32'h    FFF00393    ;    //    addi x7 x0 -1      ====        li t2, 0xffffffff
                                                  30'd    607    : data = 32'h    FFF00593    ;    //    addi x11 x0 -1      ====        li a1, 0xffffffff
                                                  30'd    608    : data = 32'h    00000813    ;    //    addi x16 x0 0      ====        li a6, 0x0
                                                  30'd    609    : data = 32'h    00000093    ;    //    addi x1 x0 0      ====        li ra, 0x0
                                                  30'd    610    : data = 32'h    00000493    ;    //    addi x9 x0 0      ====        li s1, 0x0
                                                  30'd    611    : data = 32'h    00000413    ;    //    addi x8 x0 0      ====        li s0, 0x0
                                                  30'd    612    : data = 32'h    5A8F3697    ;    //    auipc x13 370931      ====        auipc a3, 370931
                                                  30'd    613    : data = 32'h    52793617    ;    //    auipc x12 337811      ====        auipc a2, 337811
                                                  30'd    614    : data = 32'h    6AB41097    ;    //    auipc x1 437057      ====        auipc ra, 437057
                                                  30'd    615    : data = 32'h    30D60913    ;    //    addi x18 x12 781      ====        addi s2, a2, 781
                                                  30'd    616    : data = 32'h    008586B3    ;    //    add x13 x11 x8      ====        add a3, a1, s0
                                                  30'd    617    : data = 32'h    FC160913    ;    //    addi x18 x12 -63      ====        addi s2, a2, -63
                                                  30'd    618    : data = 32'h    BBBD3837    ;    //    lui x16 768979      ====        lui a6, 768979
                                                  30'd    619    : data = 32'h    E24E3937    ;    //    lui x18 926947      ====        lui s2, 926947
                                                  30'd    620    : data = 32'h    64E0A5B7    ;    //    lui x11 413194      ====        lui a1, 413194
                                                  30'd    621    : data = 32'h    49365837    ;    //    lui x16 299877      ====        lui a6, 299877
                                                  30'd    622    : data = 32'h    6FB58613    ;    //    addi x12 x11 1787      ====        addi a2, a1, 1787
                                                  30'd    623    : data = 32'h    26438913    ;    //    addi x18 x7 612      ====        addi s2, t2, 612
                                                  30'd    624    : data = 32'h    31C40913    ;    //    addi x18 x8 796      ====        addi s2, s0, 796
                                                  30'd    625    : data = 32'h    010080B3    ;    //    add x1 x1 x16      ====        add ra, ra, a6
                                                  30'd    626    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    627    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    628    : data = 32'h    73F90613    ;    //    addi x12 x18 1855      ====        addi a2, s2, 1855
                                                  30'd    629    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    630    : data = 32'h    1FE77397    ;    //    auipc x7 130679      ====        auipc t2, 130679
                                                //  30'd    631    : data = 32'h    50D0A0EF    ;    //    jal x1 44300      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_20
                                                  30'd    632    : data = 32'h    437B88B7    ;    //    lui x17 276408      ====        li a7, 0x437b781e #start riscv_int_numeric_corner_stream_25
                                                  30'd    633    : data = 32'h    81E88893    ;    //    addi x17 x17 -2018      ====        li a7, 0x437b781e #start riscv_int_numeric_corner_stream_25
                                                  30'd    634    : data = 32'h    FFF00313    ;    //    addi x6 x0 -1      ====        li t1, 0xffffffff
                                                  30'd    635    : data = 32'h    FFF00E93    ;    //    addi x29 x0 -1      ====        li t4, 0xffffffff
                                                  30'd    636    : data = 32'h    2E887E37    ;    //    lui x28 190599      ====        li t3, 0x2e8870b3
                                                  30'd    637    : data = 32'h    0B3E0E13    ;    //    addi x28 x28 179      ====        li t3, 0x2e8870b3
                                                  30'd    638    : data = 32'h    00000493    ;    //    addi x9 x0 0      ====        li s1, 0x0
                                                  30'd    639    : data = 32'h    FFF00613    ;    //    addi x12 x0 -1      ====        li a2, 0xffffffff
                                                  30'd    640    : data = 32'h    FFF00F93    ;    //    addi x31 x0 -1      ====        li t6, 0xffffffff
                                                  30'd    641    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff
                                                  30'd    642    : data = 32'h    FFF00C93    ;    //    addi x25 x0 -1      ====        li s9, 0xffffffff
                                                  30'd    643    : data = 32'h    00000D13    ;    //    addi x26 x0 0      ====        li s10, 0x0
                                                  30'd    644    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    645    : data = 32'h    01C08EB3    ;    //    add x29 x1 x28      ====        add t4, ra, t3
                                                  30'd    646    : data = 32'h    00C608B3    ;    //    add x17 x12 x12      ====        add a7, a2, a2
                                                  30'd    647    : data = 32'h    7FE40E97    ;    //    auipc x29 523840      ====        auipc t4, 523840
                                                  30'd    648    : data = 32'h    01C308B3    ;    //    add x17 x6 x28      ====        add a7, t1, t3
                                                  30'd    649    : data = 32'h    A088AD37    ;    //    lui x26 657546      ====        lui s10, 657546
                                                  30'd    650    : data = 32'h    B81E0613    ;    //    addi x12 x28 -1151      ====        addi a2, t3, -1151
                                                  30'd    651    : data = 32'h    01AD0EB3    ;    //    add x29 x26 x26      ====        add t4, s10, s10
                                                  30'd    652    : data = 32'h    F7388893    ;    //    addi x17 x17 -141      ====        addi a7, a7, -141
                                                  30'd    653    : data = 32'h    F8FEB897    ;    //    auipc x17 1019883      ====        auipc a7, 1019883
                                                  30'd    654    : data = 32'h    011880B3    ;    //    add x1 x17 x17      ====        add ra, a7, a7
                                                  30'd    655    : data = 32'h    06E30093    ;    //    addi x1 x6 110      ====        addi ra, t1, 110
                                                  30'd    656    : data = 32'h    0FFE8E13    ;    //    addi x28 x29 255      ====        addi t3, t4, 255
                                                  30'd    657    : data = 32'h    10871097    ;    //    auipc x1 67697      ====        auipc ra, 67697
                                                  30'd    658    : data = 32'h    01A30E33    ;    //    add x28 x6 x26      ====        add t3, t1, s10
                                                  30'd    659    : data = 32'h    009F8633    ;    //    add x12 x31 x9      ====        add a2, t6, s1
                                                  30'd    660    : data = 32'h    73298FB7    ;    //    lui x31 471704      ====        lui t6, 471704
                                                  30'd    661    : data = 32'h    09C48F93    ;    //    addi x31 x9 156      ====        addi t6, s1, 156
                                                  30'd    662    : data = 32'h    6FFE0897    ;    //    auipc x17 458720      ====        auipc a7, 458720
                                                  30'd    663    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                 // 30'd    664    : data = 32'h    4890A0EF    ;    //    jal x1 44168      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_25
                                                  30'd    665    : data = 32'h    800008B7    ;    //    lui x17 524288      ====        li a7, 0x80000000 #start riscv_int_numeric_corner_stream_3
                                                  30'd    666    : data = 32'h    00088893    ;    //    addi x17 x17 0      ====        li a7, 0x80000000 #start riscv_int_numeric_corner_stream_3
                                                  30'd    667    : data = 32'h    FFF00B13    ;    //    addi x22 x0 -1      ====        li s6, 0xffffffff
                                                  30'd    668    : data = 32'h    80000CB7    ;    //    lui x25 524288      ====        li s9, 0x80000000
                                                  30'd    669    : data = 32'h    000C8C93    ;    //    addi x25 x25 0      ====        li s9, 0x80000000
                                                  30'd    670    : data = 32'h    FFF00613    ;    //    addi x12 x0 -1      ====        li a2, 0xffffffff
                                                  30'd    671    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff
                                                  30'd    672    : data = 32'h    FFF00813    ;    //    addi x16 x0 -1      ====        li a6, 0xffffffff
                                                  30'd    673    : data = 32'h    FFF00313    ;    //    addi x6 x0 -1      ====        li t1, 0xffffffff
                                                  30'd    674    : data = 32'h    00000493    ;    //    addi x9 x0 0      ====        li s1, 0x0
                                                  30'd    675    : data = 32'h    00000693    ;    //    addi x13 x0 0      ====        li a3, 0x0
                                                  30'd    676    : data = 32'h    FFF00B93    ;    //    addi x23 x0 -1      ====        li s7, 0xffffffff
                                                  30'd    677    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    678    : data = 32'h    D755DB97    ;    //    auipc x23 882013      ====        auipc s7, 882013
                                                  30'd    679    : data = 32'h    5C8CE337    ;    //    lui x6 379086      ====        lui t1, 379086
                                                  30'd    680    : data = 32'h    97DB8813    ;    //    addi x16 x23 -1667      ====        addi a6, s7, -1667
                                                  30'd    681    : data = 32'h    0C425497    ;    //    auipc x9 50213      ====        auipc s1, 50213
                                                  30'd    682    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    683    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    684    : data = 32'h    B55CE617    ;    //    auipc x12 742862      ====        auipc a2, 742862
                                                  30'd    685    : data = 32'h    C728F837    ;    //    lui x16 815759      ====        lui a6, 815759
                                                  30'd    686    : data = 32'h    00130CB3    ;    //    add x25 x6 x1      ====        add s9, t1, ra
                                                  30'd    687    : data = 32'h    B770CB97    ;    //    auipc x23 751372      ====        auipc s7, 751372
                                                  30'd    688    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    689    : data = 32'h    00D68BB3    ;    //    add x23 x13 x13      ====        add s7, a3, a3
                                                  30'd    690    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    691    : data = 32'h    7526CB97    ;    //    auipc x23 479852      ====        auipc s7, 479852
                                                  30'd    692    : data = 32'h    016B8CB3    ;    //    add x25 x23 x22      ====        add s9, s7, s6
                                                  30'd    693    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    694    : data = 32'h    410B8B33    ;    //    sub x22 x23 x16      ====        sub s6, s7, a6
                                                  30'd    695    : data = 32'h    1460C0B7    ;    //    lui x1 83468      ====        lui ra, 83468
                                                  30'd    696    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    697    : data = 32'h    40180833    ;    //    sub x16 x16 x1      ====        sub a6, a6, ra
                                                  30'd    698    : data = 32'h    CB9E76B7    ;    //    lui x13 834023      ====        lui a3, 834023
                                                  30'd    699    : data = 32'h    0CB34697    ;    //    auipc x13 52020      ====        auipc a3, 52020
                                                  30'd    700    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    701    : data = 32'h    0AB51B37    ;    //    lui x22 43857      ====        lui s6, 43857
                                                  30'd    702    : data = 32'h    411800B3    ;    //    sub x1 x16 x17      ====        sub ra, a6, a7
                                                  30'd    703    : data = 32'h    410808B3    ;    //    sub x17 x16 x16      ====        sub a7, a6, a6
                                                  30'd    704    : data = 32'h    00C80B33    ;    //    add x22 x16 x12      ====        add s6, a6, a2
                                                 // 30'd    705    : data = 32'h    3E50A0EF    ;    //    jal x1 44004      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_3
                                                  30'd    706    : data = 32'h    FFF00C13    ;    //    addi x24 x0 -1      ====        li s8, 0xffffffff #start riscv_int_numeric_corner_stream_35
                                                  30'd    707    : data = 32'h    00000693    ;    //    addi x13 x0 0      ====        li a3, 0x0
                                                  30'd    708    : data = 32'h    80000437    ;    //    lui x8 524288      ====        li s0, 0x80000000
                                                  30'd    709    : data = 32'h    00040413    ;    //    addi x8 x8 0      ====        li s0, 0x80000000
                                                  30'd    710    : data = 32'h    FFF00113    ;    //    addi x2 x0 -1      ====        li sp, 0xffffffff
                                                  30'd    711    : data = 32'h    00000993    ;    //    addi x19 x0 0      ====        li s3, 0x0
                                                  30'd    712    : data = 32'h    FFF00913    ;    //    addi x18 x0 -1      ====        li s2, 0xffffffff
                                                  30'd    713    : data = 32'h    83C533B7    ;    //    lui x7 539731      ====        li t2, 0x83c5299f
                                                  30'd    714    : data = 32'h    99F38393    ;    //    addi x7 x7 -1633      ====        li t2, 0x83c5299f
                                                  30'd    715    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff
                                                  30'd    716    : data = 32'h    FFF00493    ;    //    addi x9 x0 -1      ====        li s1, 0xffffffff
                                                  30'd    717    : data = 32'h    00000E13    ;    //    addi x28 x0 0      ====        li t3, 0x0
                                                  30'd    718    : data = 32'h    05FE0413    ;    //    addi x8 x28 95      ====        addi s0, t3, 95
                                                  30'd    719    : data = 32'h    40D98E33    ;    //    sub x28 x19 x13      ====        sub t3, s3, a3
                                                  30'd    720    : data = 32'h    ED364497    ;    //    auipc x9 971620      ====        auipc s1, 971620
                                                  30'd    721    : data = 32'h    B65B2417    ;    //    auipc x8 746930      ====        auipc s0, 746930
                                                  30'd    722    : data = 32'h    FA763C37    ;    //    lui x24 1025891      ====        lui s8, 1025891
                                                  30'd    723    : data = 32'h    41CE0433    ;    //    sub x8 x28 x28      ====        sub s0, t3, t3
                                                  30'd    724    : data = 32'h    402980B3    ;    //    sub x1 x19 x2      ====        sub ra, s3, sp
                                                  30'd    725    : data = 32'h    02E98693    ;    //    addi x13 x19 46      ====        addi a3, s3, 46
                                                  30'd    726    : data = 32'h    93FD2E37    ;    //    lui x28 606162      ====        lui t3, 606162
                                                  30'd    727    : data = 32'h    0B046137    ;    //    lui x2 45126      ====        lui sp, 45126
                                                  30'd    728    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    729    : data = 32'h    013983B3    ;    //    add x7 x19 x19      ====        add t2, s3, s3
                                                  30'd    730    : data = 32'h    41238C33    ;    //    sub x24 x7 x18      ====        sub s8, t2, s2
                                                  30'd    731    : data = 32'h    1C319137    ;    //    lui x2 115481      ====        lui sp, 115481
                                                  30'd    732    : data = 32'h    41238E33    ;    //    sub x28 x7 x18      ====        sub t3, t2, s2
                                                  30'd    733    : data = 32'h    A9208993    ;    //    addi x19 x1 -1390      ====        addi s3, ra, -1390
                                                  30'd    734    : data = 32'h    01CC09B3    ;    //    add x19 x24 x28      ====        add s3, s8, t3
                                                  30'd    735    : data = 32'h    1CD19E37    ;    //    lui x28 118041      ====        lui t3, 118041
                                                  30'd    736    : data = 32'h    3FC38913    ;    //    addi x18 x7 1020      ====        addi s2, t2, 1020
                                                  30'd    737    : data = 32'h    780F7E37    ;    //    lui x28 491767      ====        lui t3, 491767
                                                  30'd    738    : data = 32'h    E0298693    ;    //    addi x13 x19 -510      ====        addi a3, s3, -510
                                                  30'd    739    : data = 32'h    40248133    ;    //    sub x2 x9 x2      ====        sub sp, s1, sp
                                                  30'd    740    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    741    : data = 32'h    007983B3    ;    //    add x7 x19 x7      ====        add t2, s3, t2
                                                  30'd    742    : data = 32'h    947F1E37    ;    //    lui x28 608241      ====        lui t3, 608241
                                                  30'd    743    : data = 32'h    01290433    ;    //    add x8 x18 x18      ====        add s0, s2, s2
                                                  30'd    744    : data = 32'h    C106AE37    ;    //    lui x28 790634      ====        lui t3, 790634
                                               //   30'd    745    : data = 32'h    3450A0EF    ;    //    jal x1 43844      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_35
                                                  30'd    746    : data = 32'h    00B4C7B7    ;    //    lui x15 2892      ====        li a5, 0xb4c19b #start riscv_int_numeric_corner_stream_15
                                                  30'd    747    : data = 32'h    19B78793    ;    //    addi x15 x15 411      ====        li a5, 0xb4c19b #start riscv_int_numeric_corner_stream_15
                                                  30'd    748    : data = 32'h    80000437    ;    //    lui x8 524288      ====        li s0, 0x80000000
                                                  30'd    749    : data = 32'h    00040413    ;    //    addi x8 x8 0      ====        li s0, 0x80000000
                                                  30'd    750    : data = 32'h    00000E13    ;    //    addi x28 x0 0      ====        li t3, 0x0
                                                  30'd    751    : data = 32'h    80000737    ;    //    lui x14 524288      ====        li a4, 0x80000000
                                                  30'd    752    : data = 32'h    00070713    ;    //    addi x14 x14 0      ====        li a4, 0x80000000
                                                  30'd    753    : data = 32'h    00000093    ;    //    addi x1 x0 0      ====        li ra, 0x0
                                                  30'd    754    : data = 32'h    FFF00693    ;    //    addi x13 x0 -1      ====        li a3, 0xffffffff
                                                  30'd    755    : data = 32'h    FFF00893    ;    //    addi x17 x0 -1      ====        li a7, 0xffffffff
                                                  30'd    756    : data = 32'h    96D13AB7    ;    //    lui x21 617747      ====        li s5, 0x96d12823
                                                  30'd    757    : data = 32'h    823A8A93    ;    //    addi x21 x21 -2013      ====        li s5, 0x96d12823
                                                  30'd    758    : data = 32'h    80000CB7    ;    //    lui x25 524288      ====        li s9, 0x80000000
                                                  30'd    759    : data = 32'h    000C8C93    ;    //    addi x25 x25 0      ====        li s9, 0x80000000
                                                  30'd    760    : data = 32'h    800003B7    ;    //    lui x7 524288      ====        li t2, 0x80000000
                                                  30'd    761    : data = 32'h    00038393    ;    //    addi x7 x7 0      ====        li t2, 0x80000000
                                                  30'd    762    : data = 32'h    40F083B3    ;    //    sub x7 x1 x15      ====        sub t2, ra, a5
                                                  30'd    763    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    764    : data = 32'h    001C87B3    ;    //    add x15 x25 x1      ====        add a5, s9, ra
                                                  30'd    765    : data = 32'h    A53CB797    ;    //    auipc x15 676811      ====        auipc a5, 676811
                                                  30'd    766    : data = 32'h    58ADE437    ;    //    lui x8 363230      ====        lui s0, 363230
                                                  30'd    767    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    768    : data = 32'h    F5039AB7    ;    //    lui x21 1003577      ====        lui s5, 1003577
                                                  30'd    769    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    770    : data = 32'h    C1EC8E13    ;    //    addi x28 x25 -994      ====        addi t3, s9, -994
                                                  30'd    771    : data = 32'h    2C7716B7    ;    //    lui x13 182129      ====        lui a3, 182129
                                                  30'd    772    : data = 32'h    9F0D3C97    ;    //    auipc x25 651475      ====        auipc s9, 651475
                                                  30'd    773    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    774    : data = 32'h    00FA8733    ;    //    add x14 x21 x15      ====        add a4, s5, a5
                                                  30'd    775    : data = 32'h    A1438713    ;    //    addi x14 x7 -1516      ====        addi a4, t2, -1516
                                                  30'd    776    : data = 32'h    367F0797    ;    //    auipc x15 223216      ====        auipc a5, 223216
                                                  30'd    777    : data = 32'h    00D08733    ;    //    add x14 x1 x13      ====        add a4, ra, a3
                                                  30'd    778    : data = 32'h    5F0CCCB7    ;    //    lui x25 389324      ====        lui s9, 389324
                                                  30'd    779    : data = 32'h    F25343B7    ;    //    lui x7 992564      ====        lui t2, 992564
                                                  30'd    780    : data = 32'h    00F086B3    ;    //    add x13 x1 x15      ====        add a3, ra, a5
                                                  30'd    781    : data = 32'h    B7212437    ;    //    lui x8 750098      ====        lui s0, 750098
                                               //   30'd    782    : data = 32'h    2B10A0EF    ;    //    jal x1 43696      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_15
                                                  30'd    783    : data = 32'h    80000937    ;    //    lui x18 524288      ====        li s2, 0x80000000 #start riscv_int_numeric_corner_stream_13
                                                  30'd    784    : data = 32'h    00090913    ;    //    addi x18 x18 0      ====        li s2, 0x80000000 #start riscv_int_numeric_corner_stream_13
                                                  30'd    785    : data = 32'h    800008B7    ;    //    lui x17 524288      ====        li a7, 0x80000000
                                                  30'd    786    : data = 32'h    00088893    ;    //    addi x17 x17 0      ====        li a7, 0x80000000
                                                  30'd    787    : data = 32'h    80000CB7    ;    //    lui x25 524288      ====        li s9, 0x80000000
                                                  30'd    788    : data = 32'h    000C8C93    ;    //    addi x25 x25 0      ====        li s9, 0x80000000
                                                  30'd    789    : data = 32'h    00000C13    ;    //    addi x24 x0 0      ====        li s8, 0x0
                                                  30'd    790    : data = 32'h    00000313    ;    //    addi x6 x0 0      ====        li t1, 0x0
                                                  30'd    791    : data = 32'h    DC5AFDB7    ;    //    lui x27 902575      ====        li s11, 0xdc5af53e
                                                  30'd    792    : data = 32'h    53ED8D93    ;    //    addi x27 x27 1342      ====        li s11, 0xdc5af53e
                                                  30'd    793    : data = 32'h    00000793    ;    //    addi x15 x0 0      ====        li a5, 0x0
                                                  30'd    794    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff
                                                  30'd    795    : data = 32'h    00000F93    ;    //    addi x31 x0 0      ====        li t6, 0x0
                                                  30'd    796    : data = 32'h    6DDF0A37    ;    //    lui x20 450032      ====        li s4, 0x6ddefb74
                                                  30'd    797    : data = 32'h    B74A0A13    ;    //    addi x20 x20 -1164      ====        li s4, 0x6ddefb74
                                                  30'd    798    : data = 32'h    41BC0A33    ;    //    sub x20 x24 x27      ====        sub s4, s8, s11
                                                  30'd    799    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    800    : data = 32'h    411C07B3    ;    //    sub x15 x24 x17      ====        sub a5, s8, a7
                                                  30'd    801    : data = 32'h    01B880B3    ;    //    add x1 x17 x27      ====        add ra, a7, s11
                                                  30'd    802    : data = 32'h    E8A57C17    ;    //    auipc x24 952919      ====        auipc s8, 952919
                                                  30'd    803    : data = 32'h    5ADD3C97    ;    //    auipc x25 372179      ====        auipc s9, 372179
                                                  30'd    804    : data = 32'h    7B55C337    ;    //    lui x6 505180      ====        lui t1, 505180
                                                  30'd    805    : data = 32'h    01BD8C33    ;    //    add x24 x27 x27      ====        add s8, s11, s11
                                                  30'd    806    : data = 32'h    931D2C17    ;    //    auipc x24 602578      ====        auipc s8, 602578
                                                  30'd    807    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    808    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    809    : data = 32'h    24434317    ;    //    auipc x6 148532      ====        auipc t1, 148532
                                                  30'd    810    : data = 32'h    AD350DB7    ;    //    lui x27 709456      ====        lui s11, 709456
                                                  30'd    811    : data = 32'h    A72C8C93    ;    //    addi x25 x25 -1422      ====        addi s9, s9, -1422
                                                  30'd    812    : data = 32'h    67CD8913    ;    //    addi x18 x27 1660      ====        addi s2, s11, 1660
                                                  30'd    813    : data = 32'h    01878CB3    ;    //    add x25 x15 x24      ====        add s9, a5, s8
                                                  30'd    814    : data = 32'h    CBC78797    ;    //    auipc x15 834680      ====        auipc a5, 834680
                                                  30'd    815    : data = 32'h    018880B3    ;    //    add x1 x17 x24      ====        add ra, a7, s8
                                                  30'd    816    : data = 32'h    B6BA2CB7    ;    //    lui x25 748450      ====        lui s9, 748450
			 	 default: data = 32'h00000013; 
 		endcase

	assign irdata_o = ird_i ? data : 32'h0;
	
	
endmodule
