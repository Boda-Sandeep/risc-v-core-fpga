module instruction_memory (
	input  			clk_i,
	input  			reset_i,
	input  [31:0]	iaddr_i,
	input  			ird_i,
	output accept,
	output [31:0]	irdata_o
);

	reg [31:0] data; 
	assign accept =1;

	always @(posedge clk_i)
		case (iaddr_i[31:2])
		                                      //    Mem Addr      //32'h       MachineCode  ;    //	BasicCode	     ====    OriginalCode

                                                  30'd	  0	   : data = 32'h	00000013	;    //	addi x0 x0 0	  ====    	nop
                                                  30'd    1    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4    : data = 32'h    00011137     ;    // 0x0	0x00011137	lui x2 17	li, sp, 68000
                                                  30'd    5    : data = 32'h    9A010113     ;    // 0x4	0x9A010113	addi x2 x2 -1632	li, sp, 68000
                                                  30'd    6    : data = 32'h    FE010113     ;    // 0x8	0xFE010113	addi x2 x2 -32	addi sp,sp,-32
                                                  30'd    7    : data = 32'h    00812E23     ;    // 0xc	0x00812E23	sw x8 28(x2)	sw s0,28(sp)
                                                  30'd    8    : data = 32'h    02010413     ;    // 0x10	0x02010413	addi x8 x2 32	addi s0,sp,32
                                                  30'd    9    : data = 32'h    00A00793     ;    // 0x14	0x00A00793	addi x15 x0 10	li a5,10
                                                  30'd    10    : data = 32'h    FEF42623     ;    // 0x18	0xFEF42623	sw x15 -20(x8)	sw a5,-20(s0)
                                                  30'd    11    : data = 32'h    00300793     ;    // 0x1c	0x00300793	addi x15 x0 3	li a5,3
                                                  30'd    12    : data = 32'h    FEF42423     ;    // 0x20	0xFEF42423	sw x15 -24(x8)	sw a5,-24(s0)
                                                  30'd    13    : data = 32'h    FEC42703     ;    // 0x24	0xFEC42703	lw x14 -20(x8)	lw a4,-20(s0)
                                                  30'd    14    : data = 32'h    FE842783     ;    // 0x28	0xFE842783	lw x15 -24(x8)	lw a5,-24(s0)
                                                  30'd    15    : data = 32'h    00F707B3     ;    // 0x2c	0x00F707B3	add x15 x14 x15	add a5,a4,a5
                                                  30'd    16    : data = 32'h    FEF42223     ;    // 0x30	0xFEF42223	sw x15 -28(x8)	sw a5,-28(s0)
                                                  30'd    17    : data = 32'h    00000013     ;    // 0x34	0x00000013	addi x0 x0 0	nop
                                                  30'd    18    : data = 32'h    00000013     ;    // 0x38	0x00000013	addi x0 x0 0	nop
                                                  30'd    19    : data = 32'h    00000013     ;    // 0x3c	0x00000013	addi x0 x0 0	nop
                                                  30'd    20    : data = 32'h    00000013     ;    // 0x40	0x00000013	addi x0 x0 0	nop
                                                  30'd    21    : data = 32'h    00000013     ;    // 0x44	0x00000013	addi x0 x0 0	nop
                                                  30'd    22    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    23    : data = 32'h    88888437    ;    //    lui x8 559240      ====        lui x8, 0x88888
                                                  30'd    24    : data = 32'h    0080A223    ;    //    sw x8 4(x1)      ====        sw x8, 4(x1)
                                                  30'd    25    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    26    : data = 32'h    999904B7    ;    //    lui x9 629136      ====        lui x9, 0x99990
                                                  30'd    27    : data = 32'h    0090A223    ;    //    sw x9 4(x1)      ====        sw x9, 4(x1)
                                                  30'd    28    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    29    : data = 32'h    000100B7    ;    //    lui x1 16      ====        lui x1, 0x00010
                                                  30'd    30    : data = 32'h    40008093    ;    //    addi x1 x1 1024      ====        addi x1, x1, 1024
                                                  30'd    31    : data = 32'h    0040A503    ;    //    lw x10 4(x1)      ====        lw x10, 4(x1)
                                                  30'd    32    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    33    : data = 32'h    0040A583    ;    //    lw x11 4(x1)      ====        lw x11, 4(x1)
                                                  30'd    34    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    35    : data = 32'h    0040A603    ;    //    lw x12 4(x1)      ====        lw x12, 4(x1)
                                                  30'd    36    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    37    : data = 32'h    0040A683    ;    //    lw x13 4(x1)      ====        lw x13, 4(x1)
                                                  30'd    38    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    39    : data = 32'h    0040A703    ;    //    lw x14 4(x1)      ====        lw x14, 4(x1)
                                                  30'd    40    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    41    : data = 32'h    0040A783    ;    //    lw x15 4(x1)      ====        lw x15, 4(x1)
                                                  30'd    42    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    43    : data = 32'h    0040A803    ;    //    lw x16 4(x1)      ====        lw x16, 4(x1)
                                                  30'd    44    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    45    : data = 32'h    0040A883    ;    //    lw x17 4(x1)      ====        lw x17, 4(x1)
                                                  30'd    46    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                                                  30'd    47    : data = 32'h    000100B7    ;    //    lui x1 16      ====        lui x1,0x00010
                                                  30'd    48    : data = 32'h    40008093    ;    //    addi x1 x1 1024      ====        addi x1, x1, 1024
                                                  30'd    49    : data = 32'h    04008213    ;    //    addi x4 x1 64      ====        addi x4, x1, 64
                                                  30'd    50    : data = 32'h    0040A023    ;    //    sw x4 0(x1)      ====        sw x4, 0x0(x1)
                                                  30'd    51    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    52    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    53    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    54    : data = 32'h    F9A4E037    ;    //    lui x0 1022542      ====        li x0, 0xf9a4dc93
                                                  30'd    55    : data = 32'h    C9300013    ;    //    addi x0 x0 -877      ====        li x0, 0xf9a4dc93
                                                  30'd    56    : data = 32'h    27DEC0B7    ;    //    lui x1 163308      ====        li x1, 0x27debf5f
                                                  30'd    57    : data = 32'h    F5F08093    ;    //    addi x1 x1 -161      ====        li x1, 0x27debf5f
                                                  30'd    58    : data = 32'h    00F00113    ;    //    addi x2 x0 15      ====        li x2, 0xf
                                                  30'd    59    : data = 32'h    800001B7    ;    //    lui x3 524288      ====        li x3, 0x80000000
                                                  30'd    60    : data = 32'h    00018193    ;    //    addi x3 x3 0      ====        li x3, 0x80000000
                                                  30'd    61    : data = 32'h    F499D2B7    ;    //    lui x5 1001885      ====        li x5, 0xf499cae9
                                                  30'd    62    : data = 32'h    AE928293    ;    //    addi x5 x5 -1303      ====        li x5, 0xf499cae9
                                                  30'd    63    : data = 32'h    5D4DA337    ;    //    lui x6 382170      ====        li x6, 0x5d4da3ca
                                                  30'd    64    : data = 32'h    3CA30313    ;    //    addi x6 x6 970      ====        li x6, 0x5d4da3ca
                                                  30'd    65    : data = 32'h    CD62F3B7    ;    //    lui x7 841263      ====        li x7, 0xcd62ecaa
                                                  30'd    66    : data = 32'h    CAA38393    ;    //    addi x7 x7 -854      ====        li x7, 0xcd62ecaa
                                                  30'd    67    : data = 32'h    F4DD0437    ;    //    lui x8 1002960      ====        li x8, 0xf4dd0029
                                                  30'd    68    : data = 32'h    02940413    ;    //    addi x8 x8 41      ====        li x8, 0xf4dd0029
                                                  30'd    69    : data = 32'h    00C00493    ;    //    addi x9 x0 12      ====        li x9, 0xc
                                                  30'd    70    : data = 32'h    F82F4537    ;    //    lui x10 1016564      ====        li x10, 0xf82f3f90
                                                  30'd    71    : data = 32'h    F9050513    ;    //    addi x10 x10 -112      ====        li x10, 0xf82f3f90
                                                  30'd    72    : data = 32'h    B81585B7    ;    //    lui x11 754008      ====        li x11, 0xb8158480
                                                  30'd    73    : data = 32'h    48058593    ;    //    addi x11 x11 1152      ====        li x11, 0xb8158480
                                                  30'd    74    : data = 32'h    AE889637    ;    //    lui x12 714889      ====        li x12, 0xae88946d
                                                  30'd    75    : data = 32'h    46D60613    ;    //    addi x12 x12 1133      ====        li x12, 0xae88946d
                                                  30'd    76    : data = 32'h    00A00693    ;    //    addi x13 x0 10      ====        li x13, 0xa
                                                  30'd    77    : data = 32'h    00000713    ;    //    addi x14 x0 0      ====        li x14, 0x0
                                                  30'd    78    : data = 32'h    00300793    ;    //    addi x15 x0 3      ====        li x15, 0x3
                                                  30'd    79    : data = 32'h    80000837    ;    //    lui x16 524288      ====        li x16, 0x80000000
                                                  30'd    80    : data = 32'h    00080813    ;    //    addi x16 x16 0      ====        li x16, 0x80000000
                                                  30'd    81    : data = 32'h    00000893    ;    //    addi x17 x0 0      ====        li x17, 0x0
                                                  30'd    82    : data = 32'h    80000937    ;    //    lui x18 524288      ====        li x18, 0x80000000
                                                  30'd    83    : data = 32'h    00090913    ;    //    addi x18 x18 0      ====        li x18, 0x80000000
                                                  30'd    84    : data = 32'h    00B00993    ;    //    addi x19 x0 11      ====        li x19, 0xb
                                                  30'd    85    : data = 32'h    F413DA37    ;    //    lui x20 999741      ====        li x20, 0xf413c908
                                                  30'd    86    : data = 32'h    908A0A13    ;    //    addi x20 x20 -1784      ====        li x20, 0xf413c908
                                                  30'd    87    : data = 32'h    0DFF5AB7    ;    //    lui x21 57333      ====        li x21, 0xdff511b
                                                  30'd    88    : data = 32'h    11BA8A93    ;    //    addi x21 x21 283      ====        li x21, 0xdff511b
                                                  30'd    89    : data = 32'h    00000B13    ;    //    addi x22 x0 0      ====        li x22, 0x0
                                                  30'd    90    : data = 32'h    80000BB7    ;    //    lui x23 524288      ====        li x23, 0x80000000
                                                  30'd    91    : data = 32'h    000B8B93    ;    //    addi x23 x23 0      ====        li x23, 0x80000000
                                                  30'd    92    : data = 32'h    FBCDDC37    ;    //    lui x24 1031389      ====        li x24, 0xfbcdd417
                                                  30'd    93    : data = 32'h    417C0C13    ;    //    addi x24 x24 1047      ====        li x24, 0xfbcdd417
                                                  30'd    94    : data = 32'h    00000C93    ;    //    addi x25 x0 0      ====        li x25, 0x0
                                                  30'd    95    : data = 32'h    91240D37    ;    //    lui x26 594496      ====        li x26, 0x9123f832
                                                  30'd    96    : data = 32'h    832D0D13    ;    //    addi x26 x26 -1998      ====        li x26, 0x9123f832
                                                  30'd    97    : data = 32'h    80000DB7    ;    //    lui x27 524288      ====        li x27, 0x80000000
                                                  30'd    98    : data = 32'h    000D8D93    ;    //    addi x27 x27 0      ====        li x27, 0x80000000
                                                  30'd    99    : data = 32'h    80000E37    ;    //    lui x28 524288      ====        li x28, 0x80000000
                                                  30'd    100    : data = 32'h    000E0E13    ;    //    addi x28 x28 0      ====        li x28, 0x80000000
                                                  30'd    101    : data = 32'h    80000EB7    ;    //    lui x29 524288      ====        li x29, 0x80000000
                                                  30'd    102    : data = 32'h    000E8E93    ;    //    addi x29 x29 0      ====        li x29, 0x80000000
                                                  30'd    103    : data = 32'h    1AD0CFB7    ;    //    lui x31 109836      ====        li x31, 0x1ad0bd45
                                                  30'd    104    : data = 32'h    D45F8F93    ;    //    addi x31 x31 -699      ====        li x31, 0x1ad0bd45
                                                  30'd    105    : data = 32'h    800007B7    ;    //    lui x15 524288      ====        main: li a5, 0x80000000 #start riscv_int_numeric_corner_stream_10
                                                  30'd    106    : data = 32'h    00078793    ;    //    addi x15 x15 0      ====        main: li a5, 0x80000000 #start riscv_int_numeric_corner_stream_10
                                                  30'd    107    : data = 32'h    5A10D937    ;    //    lui x18 368909      ====        li s2, 0x5a10d661
                                                  30'd    108    : data = 32'h    66190913    ;    //    addi x18 x18 1633      ====        li s2, 0x5a10d661
                                                  30'd    109    : data = 32'h    FFF00413    ;    //    addi x8 x0 -1      ====        li s0, 0xffffffff
                                                  30'd    110    : data = 32'h    00000E93    ;    //    addi x29 x0 0      ====        li t4, 0x0
                                                  30'd    111    : data = 32'h    FFF00893    ;    //    addi x17 x0 -1      ====        li a7, 0xffffffff
                                                  30'd    112    : data = 32'h    35049CB7    ;    //    lui x25 217161      ====        li s9, 0x35049129
                                                  30'd    113    : data = 32'h    129C8C93    ;    //    addi x25 x25 297      ====        li s9, 0x35049129
                                                  30'd    114    : data = 32'h    FFF00393    ;    //    addi x7 x0 -1      ====        li t2, 0xffffffff
                                                  30'd    115    : data = 32'h    410546B7    ;    //    lui x13 266324      ====        li a3, 0x41053ec0
                                                  30'd    116    : data = 32'h    EC068693    ;    //    addi x13 x13 -320      ====        li a3, 0x41053ec0
                                                  30'd    117    : data = 32'h    D6124637    ;    //    lui x12 876836      ====        li a2, 0xd61247be
                                                  30'd    118    : data = 32'h    7BE60613    ;    //    addi x12 x12 1982      ====        li a2, 0xd61247be
                                                  30'd    119    : data = 32'h    BA354137    ;    //    lui x2 762708      ====        li sp, 0xba353e9c
                                                  30'd    120    : data = 32'h    E9C10113    ;    //    addi x2 x2 -356      ====        li sp, 0xba353e9c
                                                  30'd    121    : data = 32'h    01D78933    ;    //    add x18 x15 x29      ====        add s2, a5, t4
                                                  30'd    122    : data = 32'h    00C10133    ;    //    add x2 x2 x12      ====        add sp, sp, a2
                                                  30'd    123    : data = 32'h    007887B3    ;    //    add x15 x17 x7      ====        add a5, a7, t2
                                                  30'd    124    : data = 32'h    008908B3    ;    //    add x17 x18 x8      ====        add a7, s2, s0
                                                  30'd    125    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    126    : data = 32'h    412687B3    ;    //    sub x15 x13 x18      ====        sub a5, a3, s2
                                                  30'd    127    : data = 32'h    40288CB3    ;    //    sub x25 x17 x2      ====        sub s9, a7, sp
                                                  30'd    128    : data = 32'h    00F38EB3    ;    //    add x29 x7 x15      ====        add t4, t2, a5
                                                  30'd    129    : data = 32'h    8B8C8393    ;    //    addi x7 x25 -1864      ====        addi t2, s9, -1864
                                                  30'd    130    : data = 32'h    71FCDCB7    ;    //    lui x25 466893      ====        lui s9, 466893
                                                  30'd    131    : data = 32'h    61CE1E97    ;    //    auipc x29 400609      ====        auipc t4, 400609
                                                  30'd    132    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    133    : data = 32'h    4564DCB7    ;    //    lui x25 284237      ====        lui s9, 284237
                                                  30'd    134    : data = 32'h    01910EB3    ;    //    add x29 x2 x25      ====        add t4, sp, s9
                                                  30'd    135    : data = 32'h    00C90613    ;    //    addi x12 x18 12      ====        addi a2, s2, 12
                                                  30'd    136    : data = 32'h    92C4D117    ;    //    auipc x2 601165      ====        auipc sp, 601165
                                                  30'd    137    : data = 32'h    4AD40613    ;    //    addi x12 x8 1197      ====        addi a2, s0, 1197
                                                  30'd    138    : data = 32'h    40740CB3    ;    //    sub x25 x8 x7      ====        sub s9, s0, t2
                                                  30'd    139    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    140    : data = 32'h    A9E10917    ;    //    auipc x18 695824      ====        auipc s2, 695824
                                                  30'd    141    : data = 32'h    41938EB3    ;    //    sub x29 x7 x25      ====        sub t4, t2, s9
                                                  30'd    142    : data = 32'h    419608B3    ;    //    sub x17 x12 x25      ====        sub a7, a2, s9
                                                  30'd    143    : data = 32'h    BE888913    ;    //    addi x18 x17 -1048      ====        addi s2, a7, -1048
                                                  30'd    144    : data = 32'h    328D17B7    ;    //    lui x15 207057      ====        lui a5, 207057
                                                  30'd    145    : data = 32'h    7DD90113    ;    //    addi x2 x18 2013      ====        addi sp, s2, 2013
                                                  30'd    146    : data = 32'h    40C90633    ;    //    sub x12 x18 x12      ====        sub a2, s2, a2
                                                  30'd    147    : data = 32'h    8BF78893    ;    //    addi x17 x15 -1857      ====        addi a7, a5, -1857
                                                  30'd    148    : data = 32'h    41288EB3    ;    //    sub x29 x17 x18      ====        sub t4, a7, s2
                                                  30'd    149    : data = 32'h    0F8577B7    ;    //    lui x15 63575      ====        lui a5, 63575
                                                  30'd    150    : data = 32'h    407E87B3    ;    //    sub x15 x29 x7      ====        sub a5, t4, t2
                                                  30'd    151    : data = 32'h    48C0B0EF    ;    //    jal x1 46220      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_10
                                                  30'd    152    : data = 32'h    800007B7    ;    //    lui x15 524288      ====        li a5, 0x80000000 #start riscv_int_numeric_corner_stream_22
                                                  30'd    153    : data = 32'h    00078793    ;    //    addi x15 x15 0      ====        li a5, 0x80000000 #start riscv_int_numeric_corner_stream_22
                                                  30'd    154    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff
                                                  30'd    155    : data = 32'h    FFF00293    ;    //    addi x5 x0 -1      ====        li t0, 0xffffffff
                                                  30'd    156    : data = 32'h    80000DB7    ;    //    lui x27 524288      ====        li s11, 0x80000000
                                                  30'd    157    : data = 32'h    000D8D93    ;    //    addi x27 x27 0      ====        li s11, 0x80000000
                                                  30'd    158    : data = 32'h    157C1A37    ;    //    lui x20 88001      ====        li s4, 0x157c126d
                                                  30'd    159    : data = 32'h    26DA0A13    ;    //    addi x20 x20 621      ====        li s4, 0x157c126d
                                                  30'd    160    : data = 32'h    80000D37    ;    //    lui x26 524288      ====        li s10, 0x80000000
                                                  30'd    161    : data = 32'h    000D0D13    ;    //    addi x26 x26 0      ====        li s10, 0x80000000
                                                  30'd    162    : data = 32'h    00000C13    ;    //    addi x24 x0 0      ====        li s8, 0x0
                                                  30'd    163    : data = 32'h    80000AB7    ;    //    lui x21 524288      ====        li s5, 0x80000000
                                                  30'd    164    : data = 32'h    000A8A93    ;    //    addi x21 x21 0      ====        li s5, 0x80000000
                                                  30'd    165    : data = 32'h    800006B7    ;    //    lui x13 524288      ====        li a3, 0x80000000
                                                  30'd    166    : data = 32'h    00068693    ;    //    addi x13 x13 0      ====        li a3, 0x80000000
                                                  30'd    167    : data = 32'h    00000193    ;    //    addi x3 x0 0      ====        li gp, 0x0
                                                  30'd    168    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    169    : data = 32'h    C2BF6D37    ;    //    lui x26 797686      ====        lui s10, 797686
                                                  30'd    170    : data = 32'h    403D06B3    ;    //    sub x13 x26 x3      ====        sub a3, s10, gp
                                                  30'd    171    : data = 32'h    1BBD0C13    ;    //    addi x24 x26 443      ====        addi s8, s10, 443
                                                  30'd    172    : data = 32'h    EF818797    ;    //    auipc x15 981016      ====        auipc a5, 981016
                                                  30'd    173    : data = 32'h    0DD28693    ;    //    addi x13 x5 221      ====        addi a3, t0, 221
                                                  30'd    174    : data = 32'h    00DD86B3    ;    //    add x13 x27 x13      ====        add a3, s11, a3
                                                  30'd    175    : data = 32'h    722D8A13    ;    //    addi x20 x27 1826      ====        addi s4, s11, 1826
                                                  30'd    176    : data = 32'h    9B00C797    ;    //    auipc x15 634892      ====        auipc a5, 634892
                                                  30'd    177    : data = 32'h    01878D33    ;    //    add x26 x15 x24      ====        add s10, a5, s8
                                                  30'd    178    : data = 32'h    CD9C0C13    ;    //    addi x24 x24 -807      ====        addi s8, s8, -807
                                                  30'd    179    : data = 32'h    9FD5B797    ;    //    auipc x15 654683      ====        auipc a5, 654683
                                                  30'd    180    : data = 32'h    5BBFC797    ;    //    auipc x15 375804      ====        auipc a5, 375804
                                                  30'd    181    : data = 32'h    F39D8D93    ;    //    addi x27 x27 -199      ====        addi s11, s11, -199
                                                  30'd    182    : data = 32'h    D24B5DB7    ;    //    lui x27 861365      ====        lui s11, 861365
                                                  30'd    183    : data = 32'h    C46A0D93    ;    //    addi x27 x20 -954      ====        addi s11, s4, -954
                                                  30'd    184    : data = 32'h    D2261AB7    ;    //    lui x21 860769      ====        lui s5, 860769
                                                  30'd    185    : data = 32'h    5C708C13    ;    //    addi x24 x1 1479      ====        addi s8, ra, 1479
                                                  30'd    186    : data = 32'h    CBB5F197    ;    //    auipc x3 834399      ====        auipc gp, 834399
                                                  30'd    187    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    188    : data = 32'h    3F80B0EF    ;    //    jal x1 46072      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_22
                                                  30'd    189    : data = 32'h    2536AC37    ;    //    lui x24 152426      ====        li s8, 0x25369e12 #start riscv_int_numeric_corner_stream_4
                                                  30'd    190    : data = 32'h    E12C0C13    ;    //    addi x24 x24 -494      ====        li s8, 0x25369e12 #start riscv_int_numeric_corner_stream_4
                                                  30'd    191    : data = 32'h    65C67EB7    ;    //    lui x29 416871      ====        li t4, 0x65c66cfd
                                                  30'd    192    : data = 32'h    CFDE8E93    ;    //    addi x29 x29 -771      ====        li t4, 0x65c66cfd
                                                  30'd    193    : data = 32'h    00000E13    ;    //    addi x28 x0 0      ====        li t3, 0x0
                                                  30'd    194    : data = 32'h    FFF00993    ;    //    addi x19 x0 -1      ====        li s3, 0xffffffff
                                                  30'd    195    : data = 32'h    19059137    ;    //    lui x2 102489      ====        li sp, 0x190590fd
                                                  30'd    196    : data = 32'h    0FD10113    ;    //    addi x2 x2 253      ====        li sp, 0x190590fd
                                                  30'd    197    : data = 32'h    FFF00D13    ;    //    addi x26 x0 -1      ====        li s10, 0xffffffff
                                                  30'd    198    : data = 32'h    00000193    ;    //    addi x3 x0 0      ====        li gp, 0x0
                                                  30'd    199    : data = 32'h    F5E1A437    ;    //    lui x8 1007130      ====        li s0, 0xf5e1a1d6
                                                  30'd    200    : data = 32'h    1D640413    ;    //    addi x8 x8 470      ====        li s0, 0xf5e1a1d6
                                                  30'd    201    : data = 32'h    FFF00913    ;    //    addi x18 x0 -1      ====        li s2, 0xffffffff
                                                  30'd    202    : data = 32'h    0155C4B7    ;    //    lui x9 5468      ====        li s1, 0x155bc11
                                                  30'd    203    : data = 32'h    C1148493    ;    //    addi x9 x9 -1007      ====        li s1, 0x155bc11
                                                  30'd    204    : data = 32'h    408C0C33    ;    //    sub x24 x24 x8      ====        sub s8, s8, s0
                                                  30'd    205    : data = 32'h    3A540193    ;    //    addi x3 x8 933      ====        addi gp, s0, 933
                                                  30'd    206    : data = 32'h    E1E6D9B7    ;    //    lui x19 925293      ====        lui s3, 925293
                                                  30'd    207    : data = 32'h    B78D0193    ;    //    addi x3 x26 -1160      ====        addi gp, s10, -1160
                                                  30'd    208    : data = 32'h    009E8EB3    ;    //    add x29 x29 x9      ====        add t4, t4, s1
                                                  30'd    209    : data = 32'h    88B07137    ;    //    lui x2 559879      ====        lui sp, 559879
                                                  30'd    210    : data = 32'h    009E8933    ;    //    add x18 x29 x9      ====        add s2, t4, s1
                                                  30'd    211    : data = 32'h    41390433    ;    //    sub x8 x18 x19      ====        sub s0, s2, s3
                                                  30'd    212    : data = 32'h    F8CBD117    ;    //    auipc x2 1019069      ====        auipc sp, 1019069
                                                  30'd    213    : data = 32'h    41C18D33    ;    //    sub x26 x3 x28      ====        sub s10, gp, t3
                                                  30'd    214    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    215    : data = 32'h    00390133    ;    //    add x2 x18 x3      ====        add sp, s2, gp
                                                  30'd    216    : data = 32'h    FD018993    ;    //    addi x19 x3 -48      ====        addi s3, gp, -48
                                                  30'd    217    : data = 32'h    40840EB3    ;    //    sub x29 x8 x8      ====        sub t4, s0, s0
                                                  30'd    218    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    219    : data = 32'h    002E0E33    ;    //    add x28 x28 x2      ====        add t3, t3, sp
                                                  30'd    220    : data = 32'h    BD3D0D13    ;    //    addi x26 x26 -1069      ====        addi s10, s10, -1069
                                                  30'd    221    : data = 32'h    00840EB3    ;    //    add x29 x8 x8      ====        add t4, s0, s0
                                                  30'd    222    : data = 32'h    AB3E9C17    ;    //    auipc x24 701417      ====        auipc s8, 701417
                                                  30'd    223    : data = 32'h    37E51137    ;    //    lui x2 228945      ====        lui sp, 228945
                                                  30'd    224    : data = 32'h    A21AD937    ;    //    lui x18 663981      ====        lui s2, 663981
                                                  30'd    225    : data = 32'h    9DA24E17    ;    //    auipc x28 645668      ====        auipc t3, 645668
                                                  30'd    226    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    227    : data = 32'h    C99D7497    ;    //    auipc x9 825815      ====        auipc s1, 825815
                                                  30'd    228    : data = 32'h    1F740993    ;    //    addi x19 x8 503      ====        addi s3, s0, 503
                                                  30'd    229    : data = 32'h    91AB7137    ;    //    lui x2 596663      ====        lui sp, 596663
                                                  30'd    230    : data = 32'h    BCDC09B7    ;    //    lui x19 773568      ====        lui s3, 773568
                                                  30'd    231    : data = 32'h    95A98E13    ;    //    addi x28 x19 -1702      ====        addi t3, s3, -1702
                                                  30'd    232    : data = 32'h    3480B0EF    ;    //    jal x1 45896      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_4
                                                  30'd    233    : data = 32'h    57B5DA37    ;    //    lui x20 359261      ====        li s4, 0x57b5c8c8 #start riscv_int_numeric_corner_stream_21
                                                  30'd    234    : data = 32'h    8C8A0A13    ;    //    addi x20 x20 -1848      ====        li s4, 0x57b5c8c8 #start riscv_int_numeric_corner_stream_21
                                                  30'd    235    : data = 32'h    800006B7    ;    //    lui x13 524288      ====        li a3, 0x80000000
                                                  30'd    236    : data = 32'h    00068693    ;    //    addi x13 x13 0      ====        li a3, 0x80000000
                                                  30'd    237    : data = 32'h    49E709B7    ;    //    lui x19 302704      ====        li s3, 0x49e6fb3e
                                                  30'd    238    : data = 32'h    B3E98993    ;    //    addi x19 x19 -1218      ====        li s3, 0x49e6fb3e
                                                  30'd    239    : data = 32'h    800001B7    ;    //    lui x3 524288      ====        li gp, 0x80000000
                                                  30'd    240    : data = 32'h    00018193    ;    //    addi x3 x3 0      ====        li gp, 0x80000000
                                                  30'd    241    : data = 32'h    FB4A5637    ;    //    lui x12 1029285      ====        li a2, 0xfb4a53f9
                                                  30'd    242    : data = 32'h    3F960613    ;    //    addi x12 x12 1017      ====        li a2, 0xfb4a53f9
                                                  30'd    243    : data = 32'h    80000CB7    ;    //    lui x25 524288      ====        li s9, 0x80000000
                                                  30'd    244    : data = 32'h    000C8C93    ;    //    addi x25 x25 0      ====        li s9, 0x80000000
                                                  30'd    245    : data = 32'h    FFF00A93    ;    //    addi x21 x0 -1      ====        li s5, 0xffffffff
                                                  30'd    246    : data = 32'h    FFF00F93    ;    //    addi x31 x0 -1      ====        li t6, 0xffffffff
                                                  30'd    247    : data = 32'h    80000E37    ;    //    lui x28 524288      ====        li t3, 0x80000000
                                                  30'd    248    : data = 32'h    000E0E13    ;    //    addi x28 x28 0      ====        li t3, 0x80000000
                                                  30'd    249    : data = 32'h    FFF00913    ;    //    addi x18 x0 -1      ====        li s2, 0xffffffff
                                                  30'd    250    : data = 32'h    419F8CB3    ;    //    sub x25 x31 x25      ====        sub s9, t6, s9
                                                  30'd    251    : data = 32'h    40DE01B3    ;    //    sub x3 x28 x13      ====        sub gp, t3, a3
                                                  30'd    252    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    253    : data = 32'h    00318CB3    ;    //    add x25 x3 x3      ====        add s9, gp, gp
                                                  30'd    254    : data = 32'h    A29B6697    ;    //    auipc x13 666038      ====        auipc a3, 666038
                                                  30'd    255    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    256    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    257    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    258    : data = 32'h    0279FC97    ;    //    auipc x25 10143      ====        auipc s9, 10143
                                                  30'd    259    : data = 32'h    59B12A97    ;    //    auipc x21 367378      ====        auipc s5, 367378
                                                  30'd    260    : data = 32'h    98494E37    ;    //    lui x28 623764      ====        lui t3, 623764
                                                  30'd    261    : data = 32'h    01F68933    ;    //    add x18 x13 x31      ====        add s2, a3, t6
                                                  30'd    262    : data = 32'h    415A8CB3    ;    //    sub x25 x21 x21      ====        sub s9, s5, s5
                                                  30'd    263    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    264    : data = 32'h    015981B3    ;    //    add x3 x19 x21      ====        add gp, s3, s5
                                                  30'd    265    : data = 32'h    40390A33    ;    //    sub x20 x18 x3      ====        sub s4, s2, gp
                                                  30'd    266    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    267    : data = 32'h    D1018693    ;    //    addi x13 x3 -752      ====        addi a3, gp, -752
                                                  30'd    268    : data = 32'h    C4990A93    ;    //    addi x21 x18 -951      ====        addi s5, s2, -951
                                                  30'd    269    : data = 32'h    212FF617    ;    //    auipc x12 135935      ====        auipc a2, 135935
                                                  30'd    270    : data = 32'h    A154B937    ;    //    lui x18 660811      ====        lui s2, 660811
                                                  30'd    271    : data = 32'h    2AC0B0EF    ;    //    jal x1 45740      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_21
                                                  30'd    272    : data = 32'h    80000137    ;    //    lui x2 524288      ====        li sp, 0x80000000 #start riscv_int_numeric_corner_stream_29
                                                  30'd    273    : data = 32'h    00010113    ;    //    addi x2 x2 0      ====        li sp, 0x80000000 #start riscv_int_numeric_corner_stream_29
                                                  30'd    274    : data = 32'h    7BD0BBB7    ;    //    lui x23 507147      ====        li s7, 0x7bd0acfa
                                                  30'd    275    : data = 32'h    CFAB8B93    ;    //    addi x23 x23 -774      ====        li s7, 0x7bd0acfa
                                                  30'd    276    : data = 32'h    AF8E7CB7    ;    //    lui x25 719079      ====        li s9, 0xaf8e6f96
                                                  30'd    277    : data = 32'h    F96C8C93    ;    //    addi x25 x25 -106      ====        li s9, 0xaf8e6f96
                                                  30'd    278    : data = 32'h    FFF00593    ;    //    addi x11 x0 -1      ====        li a1, 0xffffffff
                                                  30'd    279    : data = 32'h    519FC4B7    ;    //    lui x9 334332      ====        li s1, 0x519fc133
                                                  30'd    280    : data = 32'h    13348493    ;    //    addi x9 x9 307      ====        li s1, 0x519fc133
                                                  30'd    281    : data = 32'h    80000837    ;    //    lui x16 524288      ====        li a6, 0x80000000
                                                  30'd    282    : data = 32'h    00080813    ;    //    addi x16 x16 0      ====        li a6, 0x80000000
                                                  30'd    283    : data = 32'h    F30058B7    ;    //    lui x17 995333      ====        li a7, 0xf300533f
                                                  30'd    284    : data = 32'h    33F88893    ;    //    addi x17 x17 831      ====        li a7, 0xf300533f
                                                  30'd    285    : data = 32'h    00000B13    ;    //    addi x22 x0 0      ====        li s6, 0x0
                                                  30'd    286    : data = 32'h    FFF00293    ;    //    addi x5 x0 -1      ====        li t0, 0xffffffff
                                                  30'd    287    : data = 32'h    FFF00A93    ;    //    addi x21 x0 -1      ====        li s5, 0xffffffff
                                                  30'd    288    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    289    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    290    : data = 32'h    DD080813    ;    //    addi x16 x16 -560      ====        addi a6, a6, -560
                                                  30'd    291    : data = 32'h    FE8574B7    ;    //    lui x9 1042519      ====        lui s1, 1042519
                                                  30'd    292    : data = 32'h    41780B33    ;    //    sub x22 x16 x23      ====        sub s6, a6, s7
                                                  30'd    293    : data = 32'h    010B02B3    ;    //    add x5 x22 x16      ====        add t0, s6, a6
                                                  30'd    294    : data = 32'h    40928133    ;    //    sub x2 x5 x9      ====        sub sp, t0, s1
                                                  30'd    295    : data = 32'h    B1F3FC97    ;    //    auipc x25 728895      ====        auipc s9, 728895
                                                  30'd    296    : data = 32'h    70D472B7    ;    //    lui x5 462151      ====        lui t0, 462151
                                                  30'd    297    : data = 32'h    AA428B93    ;    //    addi x23 x5 -1372      ====        addi s7, t0, -1372
                                                  30'd    298    : data = 32'h    CE258B93    ;    //    addi x23 x11 -798      ====        addi s7, a1, -798
                                                  30'd    299    : data = 32'h    B993D297    ;    //    auipc x5 760125      ====        auipc t0, 760125
                                                  30'd    300    : data = 32'h    409B02B3    ;    //    sub x5 x22 x9      ====        sub t0, s6, s1
                                                  30'd    301    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    302    : data = 32'h    11A58593    ;    //    addi x11 x11 282      ====        addi a1, a1, 282
                                                  30'd    303    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    304    : data = 32'h    010B0133    ;    //    add x2 x22 x16      ====        add sp, s6, a6
                                                  30'd    305    : data = 32'h    BA5A8813    ;    //    addi x16 x21 -1115      ====        addi a6, s5, -1115
                                                  30'd    306    : data = 32'h    40258133    ;    //    sub x2 x11 x2      ====        sub sp, a1, sp
                                                  30'd    307    : data = 32'h    01980BB3    ;    //    add x23 x16 x25      ====        add s7, a6, s9
                                                  30'd    308    : data = 32'h    40B805B3    ;    //    sub x11 x16 x11      ====        sub a1, a6, a1
                                                  30'd    309    : data = 32'h    CD242297    ;    //    auipc x5 840258      ====        auipc t0, 840258
                                                  30'd    310    : data = 32'h    2100B0EF    ;    //    jal x1 45584      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_29
                                                  30'd    311    : data = 32'h    F84CB937    ;    //    lui x18 1017035      ====        li s2, 0xf84cb455 #start riscv_int_numeric_corner_stream_37
                                                  30'd    312    : data = 32'h    45590913    ;    //    addi x18 x18 1109      ====        li s2, 0xf84cb455 #start riscv_int_numeric_corner_stream_37
                                                  30'd    313    : data = 32'h    00000B93    ;    //    addi x23 x0 0      ====        li s7, 0x0
                                                  30'd    314    : data = 32'h    12EFF2B7    ;    //    lui x5 77567      ====        li t0, 0x12efedab
                                                  30'd    315    : data = 32'h    DAB28293    ;    //    addi x5 x5 -597      ====        li t0, 0x12efedab
                                                  30'd    316    : data = 32'h    0D01A4B7    ;    //    lui x9 53274      ====        li s1, 0xd01a71b
                                                  30'd    317    : data = 32'h    71B48493    ;    //    addi x9 x9 1819      ====        li s1, 0xd01a71b
                                                  30'd    318    : data = 32'h    BC994D37    ;    //    lui x26 772500      ====        li s10, 0xbc993d4f
                                                  30'd    319    : data = 32'h    D4FD0D13    ;    //    addi x26 x26 -689      ====        li s10, 0xbc993d4f
                                                  30'd    320    : data = 32'h    00000713    ;    //    addi x14 x0 0      ====        li a4, 0x0
                                                  30'd    321    : data = 32'h    FFF00413    ;    //    addi x8 x0 -1      ====        li s0, 0xffffffff
                                                  30'd    322    : data = 32'h    80000A37    ;    //    lui x20 524288      ====        li s4, 0x80000000
                                                  30'd    323    : data = 32'h    000A0A13    ;    //    addi x20 x20 0      ====        li s4, 0x80000000
                                                  30'd    324    : data = 32'h    FFF00893    ;    //    addi x17 x0 -1      ====        li a7, 0xffffffff
                                                  30'd    325    : data = 32'h    5D1D73B7    ;    //    lui x7 381399      ====        li t2, 0x5d1d74a4
                                                  30'd    326    : data = 32'h    4A438393    ;    //    addi x7 x7 1188      ====        li t2, 0x5d1d74a4
                                                  30'd    327    : data = 32'h    5B237B97    ;    //    auipc x23 373303      ====        auipc s7, 373303
                                                  30'd    328    : data = 32'h    012288B3    ;    //    add x17 x5 x18      ====        add a7, t0, s2
                                                  30'd    329    : data = 32'h    40E40A33    ;    //    sub x20 x8 x14      ====        sub s4, s0, a4
                                                  30'd    330    : data = 32'h    01AD03B3    ;    //    add x7 x26 x26      ====        add t2, s10, s10
                                                  30'd    331    : data = 32'h    CC048293    ;    //    addi x5 x9 -832      ====        addi t0, s1, -832
                                                  30'd    332    : data = 32'h    6B6A2737    ;    //    lui x14 439970      ====        lui a4, 439970
                                                  30'd    333    : data = 32'h    BED70B93    ;    //    addi x23 x14 -1043      ====        addi s7, a4, -1043
                                                  30'd    334    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    335    : data = 32'h    7AF20717    ;    //    auipc x14 503584      ====        auipc a4, 503584
                                                  30'd    336    : data = 32'h    007404B3    ;    //    add x9 x8 x7      ====        add s1, s0, t2
                                                  30'd    337    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    338    : data = 32'h    0E8A0B93    ;    //    addi x23 x20 232      ====        addi s7, s4, 232
                                                  30'd    339    : data = 32'h    6AC86397    ;    //    auipc x7 437382      ====        auipc t2, 437382
                                                  30'd    340    : data = 32'h    412883B3    ;    //    sub x7 x17 x18      ====        sub t2, a7, s2
                                                  30'd    341    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    342    : data = 32'h    017404B3    ;    //    add x9 x8 x23      ====        add s1, s0, s7
                                                  30'd    343    : data = 32'h    7400C297    ;    //    auipc x5 475148      ====        auipc t0, 475148
                                                  30'd    344    : data = 32'h    40928433    ;    //    sub x8 x5 x9      ====        sub s0, t0, s1
                                                  30'd    345    : data = 32'h    4C387737    ;    //    lui x14 312199      ====        lui a4, 312199
                                                  30'd    346    : data = 32'h    786984B7    ;    //    lui x9 493208      ====        lui s1, 493208
                                                  30'd    347    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    348    : data = 32'h    0096B297    ;    //    auipc x5 2411      ====        auipc t0, 2411
                                                  30'd    349    : data = 32'h    A2712417    ;    //    auipc x8 665362      ====        auipc s0, 665362
                                                  30'd    350    : data = 32'h    1700B0EF    ;    //    jal x1 45424      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_37
                                                  30'd    351    : data = 32'h    45FA2337    ;    //    lui x6 286626      ====        li t1, 0x45fa2248 #start riscv_int_numeric_corner_stream_24
                                                  30'd    352    : data = 32'h    24830313    ;    //    addi x6 x6 584      ====        li t1, 0x45fa2248 #start riscv_int_numeric_corner_stream_24
                                                  30'd    353    : data = 32'h    80000AB7    ;    //    lui x21 524288      ====        li s5, 0x80000000
                                                  30'd    354    : data = 32'h    000A8A93    ;    //    addi x21 x21 0      ====        li s5, 0x80000000
                                                  30'd    355    : data = 32'h    00000393    ;    //    addi x7 x0 0      ====        li t2, 0x0
                                                  30'd    356    : data = 32'h    220C0937    ;    //    lui x18 139456      ====        li s2, 0x220bf84d
                                                  30'd    357    : data = 32'h    84D90913    ;    //    addi x18 x18 -1971      ====        li s2, 0x220bf84d
                                                  30'd    358    : data = 32'h    00000093    ;    //    addi x1 x0 0      ====        li ra, 0x0
                                                  30'd    359    : data = 32'h    FFF00113    ;    //    addi x2 x0 -1      ====        li sp, 0xffffffff
                                                  30'd    360    : data = 32'h    FFF00613    ;    //    addi x12 x0 -1      ====        li a2, 0xffffffff
                                                  30'd    361    : data = 32'h    E78C6EB7    ;    //    lui x29 948422      ====        li t4, 0xe78c6534
                                                  30'd    362    : data = 32'h    534E8E93    ;    //    addi x29 x29 1332      ====        li t4, 0xe78c6534
                                                  30'd    363    : data = 32'h    FE598B37    ;    //    lui x22 1041816      ====        li s6, 0xfe597c60
                                                  30'd    364    : data = 32'h    C60B0B13    ;    //    addi x22 x22 -928      ====        li s6, 0xfe597c60
                                                  30'd    365    : data = 32'h    FFF00193    ;    //    addi x3 x0 -1      ====        li gp, 0xffffffff
                                                  30'd    366    : data = 32'h    74810093    ;    //    addi x1 x2 1864      ====        addi ra, sp, 1864
                                                  30'd    367    : data = 32'h    007101B3    ;    //    add x3 x2 x7      ====        add gp, sp, t2
                                                  30'd    368    : data = 32'h    C41F9637    ;    //    lui x12 803321      ====        lui a2, 803321
                                                  30'd    369    : data = 32'h    685B0E93    ;    //    addi x29 x22 1669      ====        addi t4, s6, 1669
                                                  30'd    370    : data = 32'h    01DB0633    ;    //    add x12 x22 x29      ====        add a2, s6, t4
                                                  30'd    371    : data = 32'h    3E81E617    ;    //    auipc x12 256030      ====        auipc a2, 256030
                                                  30'd    372    : data = 32'h    006100B3    ;    //    add x1 x2 x6      ====        add ra, sp, t1
                                                  30'd    373    : data = 32'h    00760633    ;    //    add x12 x12 x7      ====        add a2, a2, t2
                                                  30'd    374    : data = 32'h    2D290913    ;    //    addi x18 x18 722      ====        addi s2, s2, 722
                                                  30'd    375    : data = 32'h    00160933    ;    //    add x18 x12 x1      ====        add s2, a2, ra
                                                  30'd    376    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    377    : data = 32'h    8A03EAB7    ;    //    lui x21 565310      ====        lui s5, 565310
                                                  30'd    378    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    379    : data = 32'h    2B4B0193    ;    //    addi x3 x22 692      ====        addi gp, s6, 692
                                                  30'd    380    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    381    : data = 32'h    002A8B33    ;    //    add x22 x21 x2      ====        add s6, s5, sp
                                                  30'd    382    : data = 32'h    01530633    ;    //    add x12 x6 x21      ====        add a2, t1, s5
                                                  30'd    383    : data = 32'h    41627E97    ;    //    auipc x29 267815      ====        auipc t4, 267815
                                                  30'd    384    : data = 32'h    B1EC8637    ;    //    lui x12 728776      ====        lui a2, 728776
                                                  30'd    385    : data = 32'h    01260933    ;    //    add x18 x12 x18      ====        add s2, a2, s2
                                                  30'd    386    : data = 32'h    1C6E8113    ;    //    addi x2 x29 454      ====        addi sp, t4, 454
                                                  30'd    387    : data = 32'h    1DC75B37    ;    //    lui x22 121973      ====        lui s6, 121973
                                                  30'd    388    : data = 32'h    36DD2937    ;    //    lui x18 224722      ====        lui s2, 224722
                                                  30'd    389    : data = 32'h    78156317    ;    //    auipc x6 491862      ====        auipc t1, 491862
                                                  30'd    390    : data = 32'h    41D30AB3    ;    //    sub x21 x6 x29      ====        sub s5, t1, t4
                                                  30'd    391    : data = 32'h    00338633    ;    //    add x12 x7 x3      ====        add a2, t2, gp
                                                  30'd    392    : data = 32'h    888B0093    ;    //    addi x1 x22 -1912      ====        addi ra, s6, -1912
                                                  30'd    393    : data = 32'h    40760B33    ;    //    sub x22 x12 x7      ====        sub s6, a2, t2
                                                  30'd    394    : data = 32'h    0C00B0EF    ;    //    jal x1 45248      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_24
                                                  30'd    395    : data = 32'h    80000EB7    ;    //    lui x29 524288      ====        li t4, 0x80000000 #start riscv_int_numeric_corner_stream_27
                                                  30'd    396    : data = 32'h    000E8E93    ;    //    addi x29 x29 0      ====        li t4, 0x80000000 #start riscv_int_numeric_corner_stream_27
                                                  30'd    397    : data = 32'h    D3F4B4B7    ;    //    lui x9 868171      ====        li s1, 0xd3f4aa26
                                                  30'd    398    : data = 32'h    A2648493    ;    //    addi x9 x9 -1498      ====        li s1, 0xd3f4aa26
                                                  30'd    399    : data = 32'h    0B6F10B7    ;    //    lui x1 46833      ====        li ra, 0xb6f12e8
                                                  30'd    400    : data = 32'h    2E808093    ;    //    addi x1 x1 744      ====        li ra, 0xb6f12e8
                                                  30'd    401    : data = 32'h    F7A553B7    ;    //    lui x7 1014357      ====        li t2, 0xf7a555ad
                                                  30'd    402    : data = 32'h    5AD38393    ;    //    addi x7 x7 1453      ====        li t2, 0xf7a555ad
                                                  30'd    403    : data = 32'h    80000CB7    ;    //    lui x25 524288      ====        li s9, 0x80000000
                                                  30'd    404    : data = 32'h    000C8C93    ;    //    addi x25 x25 0      ====        li s9, 0x80000000
                                                  30'd    405    : data = 32'h    FFF00F93    ;    //    addi x31 x0 -1      ====        li t6, 0xffffffff
                                                  30'd    406    : data = 32'h    00000593    ;    //    addi x11 x0 0      ====        li a1, 0x0
                                                  30'd    407    : data = 32'h    FFF00293    ;    //    addi x5 x0 -1      ====        li t0, 0xffffffff
                                                  30'd    408    : data = 32'h    00000713    ;    //    addi x14 x0 0      ====        li a4, 0x0
                                                  30'd    409    : data = 32'h    E991B137    ;    //    lui x2 956699      ====        li sp, 0xe991a96c
                                                  30'd    410    : data = 32'h    96C10113    ;    //    addi x2 x2 -1684      ====        li sp, 0xe991a96c
                                                  30'd    411    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    412    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    413    : data = 32'h    40710FB3    ;    //    sub x31 x2 x7      ====        sub t6, sp, t2
                                                  30'd    414    : data = 32'h    B3D5B0B7    ;    //    lui x1 736603      ====        lui ra, 736603
                                                  30'd    415    : data = 32'h    409F8733    ;    //    sub x14 x31 x9      ====        sub a4, t6, s1
                                                  30'd    416    : data = 32'h    F0E38713    ;    //    addi x14 x7 -242      ====        addi a4, t2, -242
                                                  30'd    417    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    418    : data = 32'h    40B583B3    ;    //    sub x7 x11 x11      ====        sub t2, a1, a1
                                                  30'd    419    : data = 32'h    DB110493    ;    //    addi x9 x2 -591      ====        addi s1, sp, -591
                                                  30'd    420    : data = 32'h    56228C93    ;    //    addi x25 x5 1378      ====        addi s9, t0, 1378
                                                  30'd    421    : data = 32'h    D8CA5137    ;    //    lui x2 887973      ====        lui sp, 887973
                                                  30'd    422    : data = 32'h    FF80C397    ;    //    auipc x7 1046540      ====        auipc t2, 1046540
                                                  30'd    423    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    424    : data = 32'h    00E385B3    ;    //    add x11 x7 x14      ====        add a1, t2, a4
                                                  30'd    425    : data = 32'h    C0A44737    ;    //    lui x14 789060      ====        lui a4, 789060
                                                  30'd    426    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    427    : data = 32'h    6A0B2737    ;    //    lui x14 434354      ====        lui a4, 434354
                                                  30'd    428    : data = 32'h    278800B7    ;    //    lui x1 161920      ====        lui ra, 161920
                                                  30'd    429    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    430    : data = 32'h    D9C38C93    ;    //    addi x25 x7 -612      ====        addi s9, t2, -612
                                                  30'd    431    : data = 32'h    A9EE1EB7    ;    //    lui x29 696033      ====        lui t4, 696033
                                                  30'd    432    : data = 32'h    40E10133    ;    //    sub x2 x2 x14      ====        sub sp, sp, a4
                                                  30'd    433    : data = 32'h    F7571137    ;    //    lui x2 1013105      ====        lui sp, 1013105
                                                  30'd    434    : data = 32'h    2D138F93    ;    //    addi x31 x7 721      ====        addi t6, t2, 721
                                                  30'd    435    : data = 32'h    22D64597    ;    //    auipc x11 142692      ====        auipc a1, 142692
                                                  30'd    436    : data = 32'h    0180B0EF    ;    //    jal x1 45080      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_27
                                                  30'd    437    : data = 32'h    FFF00393    ;    //    addi x7 x0 -1      ====        li t2, 0xffffffff #start riscv_int_numeric_corner_stream_39
                                                  30'd    438    : data = 32'h    38D299B7    ;    //    lui x19 232745      ====        li s3, 0x38d2979d
                                                  30'd    439    : data = 32'h    79D98993    ;    //    addi x19 x19 1949      ====        li s3, 0x38d2979d
                                                  30'd    440    : data = 32'h    00000A93    ;    //    addi x21 x0 0      ====        li s5, 0x0
                                                  30'd    441    : data = 32'h    00000593    ;    //    addi x11 x0 0      ====        li a1, 0x0
                                                  30'd    442    : data = 32'h    00000E13    ;    //    addi x28 x0 0      ====        li t3, 0x0
                                                  30'd    443    : data = 32'h    FFF00413    ;    //    addi x8 x0 -1      ====        li s0, 0xffffffff
                                                  30'd    444    : data = 32'h    80000137    ;    //    lui x2 524288      ====        li sp, 0x80000000
                                                  30'd    445    : data = 32'h    00010113    ;    //    addi x2 x2 0      ====        li sp, 0x80000000
                                                  30'd    446    : data = 32'h    00000893    ;    //    addi x17 x0 0      ====        li a7, 0x0
                                                  30'd    447    : data = 32'h    00000313    ;    //    addi x6 x0 0      ====        li t1, 0x0
                                                  30'd    448    : data = 32'h    FFF00293    ;    //    addi x5 x0 -1      ====        li t0, 0xffffffff
                                                  30'd    449    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    450    : data = 32'h    7510B9B7    ;    //    lui x19 479499      ====        lui s3, 479499
                                                  30'd    451    : data = 32'h    899EB997    ;    //    auipc x19 563691      ====        auipc s3, 563691
                                                  30'd    452    : data = 32'h    40B30433    ;    //    sub x8 x6 x11      ====        sub s0, t1, a1
                                                  30'd    453    : data = 32'h    CAB91997    ;    //    auipc x19 830353      ====        auipc s3, 830353
                                                  30'd    454    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    455    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    456    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    457    : data = 32'h    52AA1437    ;    //    lui x8 338593      ====        lui s0, 338593
                                                  30'd    458    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    459    : data = 32'h    FFCA8E13    ;    //    addi x28 x21 -4      ====        addi t3, s5, -4
                                                  30'd    460    : data = 32'h    013302B3    ;    //    add x5 x6 x19      ====        add t0, t1, s3
                                                  30'd    461    : data = 32'h    EC0E8297    ;    //    auipc x5 966888      ====        auipc t0, 966888
                                                  30'd    462    : data = 32'h    05784997    ;    //    auipc x19 22404      ====        auipc s3, 22404
                                                  30'd    463    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    464    : data = 32'h    005583B3    ;    //    add x7 x11 x5      ====        add t2, a1, t0
                                                  30'd    465    : data = 32'h    40630333    ;    //    sub x6 x6 x6      ====        sub t1, t1, t1
                                                  30'd    466    : data = 32'h    406288B3    ;    //    sub x17 x5 x6      ====        sub a7, t0, t1
                                                  30'd    467    : data = 32'h    4751B2B7    ;    //    lui x5 292123      ====        lui t0, 292123
                                                  30'd    468    : data = 32'h    AF030593    ;    //    addi x11 x6 -1296      ====        addi a1, t1, -1296
                                                  30'd    469    : data = 32'h    406E0433    ;    //    sub x8 x28 x6      ====        sub s0, t3, t1
                                                  30'd    470    : data = 32'h    413303B3    ;    //    sub x7 x6 x19      ====        sub t2, t1, s3
                                                  30'd    471    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    472    : data = 32'h    AF358593    ;    //    addi x11 x11 -1293      ====        addi a1, a1, -1293
                                                  30'd    473    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    474    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    475    : data = 32'h    007582B3    ;    //    add x5 x11 x7      ====        add t0, a1, t2
                                                  30'd    476    : data = 32'h    DC640413    ;    //    addi x8 x8 -570      ====        addi s0, s0, -570
                                                  30'd    477    : data = 32'h    7750A0EF    ;    //    jal x1 44916      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_39
                                                  30'd    478    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff #start riscv_int_numeric_corner_stream_9
                                                  30'd    479    : data = 32'h    80000137    ;    //    lui x2 524288      ====        li sp, 0x80000000
                                                  30'd    480    : data = 32'h    00010113    ;    //    addi x2 x2 0      ====        li sp, 0x80000000
                                                  30'd    481    : data = 32'h    00000C13    ;    //    addi x24 x0 0      ====        li s8, 0x0
                                                  30'd    482    : data = 32'h    FFF00A93    ;    //    addi x21 x0 -1      ====        li s5, 0xffffffff
                                                  30'd    483    : data = 32'h    80000B37    ;    //    lui x22 524288      ====        li s6, 0x80000000
                                                  30'd    484    : data = 32'h    000B0B13    ;    //    addi x22 x22 0      ====        li s6, 0x80000000
                                                  30'd    485    : data = 32'h    FFF00C93    ;    //    addi x25 x0 -1      ====        li s9, 0xffffffff
                                                  30'd    486    : data = 32'h    00000393    ;    //    addi x7 x0 0      ====        li t2, 0x0
                                                  30'd    487    : data = 32'h    FFF00B93    ;    //    addi x23 x0 -1      ====        li s7, 0xffffffff
                                                  30'd    488    : data = 32'h    80000637    ;    //    lui x12 524288      ====        li a2, 0x80000000
                                                  30'd    489    : data = 32'h    00060613    ;    //    addi x12 x12 0      ====        li a2, 0x80000000
                                                  30'd    490    : data = 32'h    55B2D5B7    ;    //    lui x11 351021      ====        li a1, 0x55b2ccfe
                                                  30'd    491    : data = 32'h    CFE58593    ;    //    addi x11 x11 -770      ====        li a1, 0x55b2ccfe
                                                  30'd    492    : data = 32'h    47BA2637    ;    //    lui x12 293794      ====        lui a2, 293794
                                                  30'd    493    : data = 32'h    E3463BB7    ;    //    lui x23 930915      ====        lui s7, 930915
                                                  30'd    494    : data = 32'h    002B0CB3    ;    //    add x25 x22 x2      ====        add s9, s6, sp
                                                  30'd    495    : data = 32'h    DC4D25B7    ;    //    lui x11 902354      ====        lui a1, 902354
                                                  30'd    496    : data = 32'h    F8C27117    ;    //    auipc x2 1018919      ====        auipc sp, 1018919
                                                  30'd    497    : data = 32'h    017385B3    ;    //    add x11 x7 x23      ====        add a1, t2, s7
                                                  30'd    498    : data = 32'h    9DA10A93    ;    //    addi x21 x2 -1574      ====        addi s5, sp, -1574
                                                  30'd    499    : data = 32'h    01960CB3    ;    //    add x25 x12 x25      ====        add s9, a2, s9
                                                  30'd    500    : data = 32'h    F2B0B0B7    ;    //    lui x1 994059      ====        lui ra, 994059
                                                  30'd    501    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    502    : data = 32'h    6D7AACB7    ;    //    lui x25 448426      ====        lui s9, 448426
                                                  30'd    503    : data = 32'h    CF938A93    ;    //    addi x21 x7 -775      ====        addi s5, t2, -775
                                                  30'd    504    : data = 32'h    419C80B3    ;    //    sub x1 x25 x25      ====        sub ra, s9, s9
                                                  30'd    505    : data = 32'h    21712397    ;    //    auipc x7 136978      ====        auipc t2, 136978
                                                  30'd    506    : data = 32'h    40C38AB3    ;    //    sub x21 x7 x12      ====        sub s5, t2, a2
                                                  30'd    507    : data = 32'h    00CB0133    ;    //    add x2 x22 x12      ====        add sp, s6, a2
                                                  30'd    508    : data = 32'h    01958633    ;    //    add x12 x11 x25      ====        add a2, a1, s9
                                                  30'd    509    : data = 32'h    86308C13    ;    //    addi x24 x1 -1949      ====        addi s8, ra, -1949
                                                  30'd    510    : data = 32'h    872B0613    ;    //    addi x12 x22 -1934      ====        addi a2, s6, -1934
                                                  30'd    511    : data = 32'h    2BB635B7    ;    //    lui x11 179043      ====        lui a1, 179043
                                                  30'd    512    : data = 32'h    33D25B37    ;    //    lui x22 212261      ====        lui s6, 212261
                                                  30'd    513    : data = 32'h    CCDE9137    ;    //    lui x2 839145      ====        lui sp, 839145
                                                  30'd    514    : data = 32'h    00BB8633    ;    //    add x12 x23 x11      ====        add a2, s7, a1
                                                  30'd    515    : data = 32'h    01658B33    ;    //    add x22 x11 x22      ====        add s6, a1, s6
                                                  30'd    516    : data = 32'h    82E6BA97    ;    //    auipc x21 536171      ====        auipc s5, 536171
                                                  30'd    517    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    518    : data = 32'h    415C8633    ;    //    sub x12 x25 x21      ====        sub a2, s9, s5
                                                  30'd    519    : data = 32'h    8520CC97    ;    //    auipc x25 545292      ====        auipc s9, 545292
                                                  30'd    520    : data = 32'h    B782C5B7    ;    //    lui x11 751660      ====        lui a1, 751660
                                                  30'd    521    : data = 32'h    6C50A0EF    ;    //    jal x1 44740      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_9
                                                  30'd    522    : data = 32'h    33525437    ;    //    lui x8 210213      ====        li s0, 0x335253fa #start riscv_int_numeric_corner_stream_26
                                                  30'd    523    : data = 32'h    3FA40413    ;    //    addi x8 x8 1018      ====        li s0, 0x335253fa #start riscv_int_numeric_corner_stream_26
                                                  30'd    524    : data = 32'h    FFF00713    ;    //    addi x14 x0 -1      ====        li a4, 0xffffffff
                                                  30'd    525    : data = 32'h    80000DB7    ;    //    lui x27 524288      ====        li s11, 0x80000000
                                                  30'd    526    : data = 32'h    000D8D93    ;    //    addi x27 x27 0      ====        li s11, 0x80000000
                                                  30'd    527    : data = 32'h    C88AF7B7    ;    //    lui x15 821423      ====        li a5, 0xc88af75b
                                                  30'd    528    : data = 32'h    75B78793    ;    //    addi x15 x15 1883      ====        li a5, 0xc88af75b
                                                  30'd    529    : data = 32'h    FFF00993    ;    //    addi x19 x0 -1      ====        li s3, 0xffffffff
                                                  30'd    530    : data = 32'h    800005B7    ;    //    lui x11 524288      ====        li a1, 0x80000000
                                                  30'd    531    : data = 32'h    00058593    ;    //    addi x11 x11 0      ====        li a1, 0x80000000
                                                  30'd    532    : data = 32'h    FFF00B93    ;    //    addi x23 x0 -1      ====        li s7, 0xffffffff
                                                  30'd    533    : data = 32'h    DDD15A37    ;    //    lui x20 908565      ====        li s4, 0xddd1523c
                                                  30'd    534    : data = 32'h    23CA0A13    ;    //    addi x20 x20 572      ====        li s4, 0xddd1523c
                                                  30'd    535    : data = 32'h    FFF00A93    ;    //    addi x21 x0 -1      ====        li s5, 0xffffffff
                                                  30'd    536    : data = 32'h    E8DF9D37    ;    //    lui x26 953849      ====        li s10, 0xe8df8e05
                                                  30'd    537    : data = 32'h    E05D0D13    ;    //    addi x26 x26 -507      ====        li s10, 0xe8df8e05
                                                  30'd    538    : data = 32'h    40BA0BB3    ;    //    sub x23 x20 x11      ====        sub s7, s4, a1
                                                  30'd    539    : data = 32'h    346B8593    ;    //    addi x11 x23 838      ====        addi a1, s7, 838
                                                  30'd    540    : data = 32'h    01AB8D33    ;    //    add x26 x23 x26      ====        add s10, s7, s10
                                                  30'd    541    : data = 32'h    103A8993    ;    //    addi x19 x21 259      ====        addi s3, s5, 259
                                                  30'd    542    : data = 32'h    A9718A17    ;    //    auipc x20 694040      ====        auipc s4, 694040
                                                  30'd    543    : data = 32'h    014A0BB3    ;    //    add x23 x20 x20      ====        add s7, s4, s4
                                                  30'd    544    : data = 32'h    40F78733    ;    //    sub x14 x15 x15      ====        sub a4, a5, a5
                                                  30'd    545    : data = 32'h    5F978D13    ;    //    addi x26 x15 1529      ====        addi s10, a5, 1529
                                                  30'd    546    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    547    : data = 32'h    CA6C4D97    ;    //    auipc x27 829124      ====        auipc s11, 829124
                                                  30'd    548    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    549    : data = 32'h    00EA0433    ;    //    add x8 x20 x14      ====        add s0, s4, a4
                                                  30'd    550    : data = 32'h    59DD5D37    ;    //    lui x26 368085      ====        lui s10, 368085
                                                  30'd    551    : data = 32'h    75A78713    ;    //    addi x14 x15 1882      ====        addi a4, a5, 1882
                                                  30'd    552    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    553    : data = 32'h    A981B5B7    ;    //    lui x11 694299      ====        lui a1, 694299
                                                  30'd    554    : data = 32'h    417B8A33    ;    //    sub x20 x23 x23      ====        sub s4, s7, s7
                                                  30'd    555    : data = 32'h    40840AB3    ;    //    sub x21 x8 x8      ====        sub s5, s0, s0
                                                  30'd    556    : data = 32'h    0C758713    ;    //    addi x14 x11 199      ====        addi a4, a1, 199
                                                  30'd    557    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    558    : data = 32'h    0D9D1417    ;    //    auipc x8 55761      ====        auipc s0, 55761
                                                  30'd    559    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    560    : data = 32'h    413D8DB3    ;    //    sub x27 x27 x19      ====        sub s11, s11, s3
                                                  30'd    561    : data = 32'h    01458433    ;    //    add x8 x11 x20      ====        add s0, a1, s4
                                                  30'd    562    : data = 32'h    F6B7DD17    ;    //    auipc x26 1010557      ====        auipc s10, 1010557
                                                  30'd    563    : data = 32'h    A0ADDD37    ;    //    lui x26 658141      ====        lui s10, 658141
                                                  30'd    564    : data = 32'h    40B98733    ;    //    sub x14 x19 x11      ====        sub a4, s3, a1
                                                  30'd    565    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    566    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    567    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    568    : data = 32'h    6090A0EF    ;    //    jal x1 44552      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_26
                                                  30'd    569    : data = 32'h    00000113    ;    //    addi x2 x0 0      ====        li sp, 0x0 #start riscv_int_numeric_corner_stream_6
                                                  30'd    570    : data = 32'h    AE9BF4B7    ;    //    lui x9 715199      ====        li s1, 0xae9bf065
                                                  30'd    571    : data = 32'h    06548493    ;    //    addi x9 x9 101      ====        li s1, 0xae9bf065
                                                  30'd    572    : data = 32'h    446D16B7    ;    //    lui x13 280273      ====        li a3, 0x446d0933
                                                  30'd    573    : data = 32'h    93368693    ;    //    addi x13 x13 -1741      ====        li a3, 0x446d0933
                                                  30'd    574    : data = 32'h    00000C93    ;    //    addi x25 x0 0      ====        li s9, 0x0
                                                  30'd    575    : data = 32'h    00000193    ;    //    addi x3 x0 0      ====        li gp, 0x0
                                                  30'd    576    : data = 32'h    FFF00B13    ;    //    addi x22 x0 -1      ====        li s6, 0xffffffff
                                                  30'd    577    : data = 32'h    B4B72FB7    ;    //    lui x31 740210      ====        li t6, 0xb4b71a5b
                                                  30'd    578    : data = 32'h    A5BF8F93    ;    //    addi x31 x31 -1445      ====        li t6, 0xb4b71a5b
                                                  30'd    579    : data = 32'h    800000B7    ;    //    lui x1 524288      ====        li ra, 0x80000000
                                                  30'd    580    : data = 32'h    00008093    ;    //    addi x1 x1 0      ====        li ra, 0x80000000
                                                  30'd    581    : data = 32'h    80000937    ;    //    lui x18 524288      ====        li s2, 0x80000000
                                                  30'd    582    : data = 32'h    00090913    ;    //    addi x18 x18 0      ====        li s2, 0x80000000
                                                  30'd    583    : data = 32'h    98D19E37    ;    //    lui x28 625945      ====        li t3, 0x98d191a8
                                                  30'd    584    : data = 32'h    1A8E0E13    ;    //    addi x28 x28 424      ====        li t3, 0x98d191a8
                                                  30'd    585    : data = 32'h    001484B3    ;    //    add x9 x9 x1      ====        add s1, s1, ra
                                                  30'd    586    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    587    : data = 32'h    3EE58B17    ;    //    auipc x22 257624      ====        auipc s6, 257624
                                                  30'd    588    : data = 32'h    A3F0BB37    ;    //    lui x22 671499      ====        lui s6, 671499
                                                  30'd    589    : data = 32'h    87CA2F97    ;    //    auipc x31 556194      ====        auipc t6, 556194
                                                  30'd    590    : data = 32'h    419E0E33    ;    //    sub x28 x28 x25      ====        sub t3, t3, s9
                                                  30'd    591    : data = 32'h    C8963F97    ;    //    auipc x31 821603      ====        auipc t6, 821603
                                                  30'd    592    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    593    : data = 32'h    33EF8E13    ;    //    addi x28 x31 830      ====        addi t3, t6, 830
                                                  30'd    594    : data = 32'h    E6555E17    ;    //    auipc x28 943445      ====        auipc t3, 943445
                                                  30'd    595    : data = 32'h    9F8ECB17    ;    //    auipc x22 653548      ====        auipc s6, 653548
                                                  30'd    596    : data = 32'h    BFC71197    ;    //    auipc x3 785521      ====        auipc gp, 785521
                                                  30'd    597    : data = 32'h    001086B3    ;    //    add x13 x1 x1      ====        add a3, ra, ra
                                                  30'd    598    : data = 32'h    97F4DE37    ;    //    lui x28 622413      ====        lui t3, 622413
                                                  30'd    599    : data = 32'h    73E68937    ;    //    lui x18 474728      ====        lui s2, 474728
                                                  30'd    600    : data = 32'h    5890A0EF    ;    //    jal x1 44424      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_6
                                                  30'd    601    : data = 32'h    00000693    ;    //    addi x13 x0 0      ====        li a3, 0x0 #start riscv_int_numeric_corner_stream_20
                                                  30'd    602    : data = 32'h    00000193    ;    //    addi x3 x0 0      ====        li gp, 0x0
                                                  30'd    603    : data = 32'h    17826637    ;    //    lui x12 96294      ====        li a2, 0x17825de0
                                                  30'd    604    : data = 32'h    DE060613    ;    //    addi x12 x12 -544      ====        li a2, 0x17825de0
                                                  30'd    605    : data = 32'h    00000913    ;    //    addi x18 x0 0      ====        li s2, 0x0
                                                  30'd    606    : data = 32'h    FFF00393    ;    //    addi x7 x0 -1      ====        li t2, 0xffffffff
                                                  30'd    607    : data = 32'h    FFF00593    ;    //    addi x11 x0 -1      ====        li a1, 0xffffffff
                                                  30'd    608    : data = 32'h    00000813    ;    //    addi x16 x0 0      ====        li a6, 0x0
                                                  30'd    609    : data = 32'h    00000093    ;    //    addi x1 x0 0      ====        li ra, 0x0
                                                  30'd    610    : data = 32'h    00000493    ;    //    addi x9 x0 0      ====        li s1, 0x0
                                                  30'd    611    : data = 32'h    00000413    ;    //    addi x8 x0 0      ====        li s0, 0x0
                                                  30'd    612    : data = 32'h    5A8F3697    ;    //    auipc x13 370931      ====        auipc a3, 370931
                                                  30'd    613    : data = 32'h    52793617    ;    //    auipc x12 337811      ====        auipc a2, 337811
                                                  30'd    614    : data = 32'h    6AB41097    ;    //    auipc x1 437057      ====        auipc ra, 437057
                                                  30'd    615    : data = 32'h    30D60913    ;    //    addi x18 x12 781      ====        addi s2, a2, 781
                                                  30'd    616    : data = 32'h    008586B3    ;    //    add x13 x11 x8      ====        add a3, a1, s0
                                                  30'd    617    : data = 32'h    FC160913    ;    //    addi x18 x12 -63      ====        addi s2, a2, -63
                                                  30'd    618    : data = 32'h    BBBD3837    ;    //    lui x16 768979      ====        lui a6, 768979
                                                  30'd    619    : data = 32'h    E24E3937    ;    //    lui x18 926947      ====        lui s2, 926947
                                                  30'd    620    : data = 32'h    64E0A5B7    ;    //    lui x11 413194      ====        lui a1, 413194
                                                  30'd    621    : data = 32'h    49365837    ;    //    lui x16 299877      ====        lui a6, 299877
                                                  30'd    622    : data = 32'h    6FB58613    ;    //    addi x12 x11 1787      ====        addi a2, a1, 1787
                                                  30'd    623    : data = 32'h    26438913    ;    //    addi x18 x7 612      ====        addi s2, t2, 612
                                                  30'd    624    : data = 32'h    31C40913    ;    //    addi x18 x8 796      ====        addi s2, s0, 796
                                                  30'd    625    : data = 32'h    010080B3    ;    //    add x1 x1 x16      ====        add ra, ra, a6
                                                  30'd    626    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    627    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    628    : data = 32'h    73F90613    ;    //    addi x12 x18 1855      ====        addi a2, s2, 1855
                                                  30'd    629    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    630    : data = 32'h    1FE77397    ;    //    auipc x7 130679      ====        auipc t2, 130679
                                                  30'd    631    : data = 32'h    50D0A0EF    ;    //    jal x1 44300      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_20
                                                  30'd    632    : data = 32'h    437B88B7    ;    //    lui x17 276408      ====        li a7, 0x437b781e #start riscv_int_numeric_corner_stream_25
                                                  30'd    633    : data = 32'h    81E88893    ;    //    addi x17 x17 -2018      ====        li a7, 0x437b781e #start riscv_int_numeric_corner_stream_25
                                                  30'd    634    : data = 32'h    FFF00313    ;    //    addi x6 x0 -1      ====        li t1, 0xffffffff
                                                  30'd    635    : data = 32'h    FFF00E93    ;    //    addi x29 x0 -1      ====        li t4, 0xffffffff
                                                  30'd    636    : data = 32'h    2E887E37    ;    //    lui x28 190599      ====        li t3, 0x2e8870b3
                                                  30'd    637    : data = 32'h    0B3E0E13    ;    //    addi x28 x28 179      ====        li t3, 0x2e8870b3
                                                  30'd    638    : data = 32'h    00000493    ;    //    addi x9 x0 0      ====        li s1, 0x0
                                                  30'd    639    : data = 32'h    FFF00613    ;    //    addi x12 x0 -1      ====        li a2, 0xffffffff
                                                  30'd    640    : data = 32'h    FFF00F93    ;    //    addi x31 x0 -1      ====        li t6, 0xffffffff
                                                  30'd    641    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff
                                                  30'd    642    : data = 32'h    FFF00C93    ;    //    addi x25 x0 -1      ====        li s9, 0xffffffff
                                                  30'd    643    : data = 32'h    00000D13    ;    //    addi x26 x0 0      ====        li s10, 0x0
                                                  30'd    644    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    645    : data = 32'h    01C08EB3    ;    //    add x29 x1 x28      ====        add t4, ra, t3
                                                  30'd    646    : data = 32'h    00C608B3    ;    //    add x17 x12 x12      ====        add a7, a2, a2
                                                  30'd    647    : data = 32'h    7FE40E97    ;    //    auipc x29 523840      ====        auipc t4, 523840
                                                  30'd    648    : data = 32'h    01C308B3    ;    //    add x17 x6 x28      ====        add a7, t1, t3
                                                  30'd    649    : data = 32'h    A088AD37    ;    //    lui x26 657546      ====        lui s10, 657546
                                                  30'd    650    : data = 32'h    B81E0613    ;    //    addi x12 x28 -1151      ====        addi a2, t3, -1151
                                                  30'd    651    : data = 32'h    01AD0EB3    ;    //    add x29 x26 x26      ====        add t4, s10, s10
                                                  30'd    652    : data = 32'h    F7388893    ;    //    addi x17 x17 -141      ====        addi a7, a7, -141
                                                  30'd    653    : data = 32'h    F8FEB897    ;    //    auipc x17 1019883      ====        auipc a7, 1019883
                                                  30'd    654    : data = 32'h    011880B3    ;    //    add x1 x17 x17      ====        add ra, a7, a7
                                                  30'd    655    : data = 32'h    06E30093    ;    //    addi x1 x6 110      ====        addi ra, t1, 110
                                                  30'd    656    : data = 32'h    0FFE8E13    ;    //    addi x28 x29 255      ====        addi t3, t4, 255
                                                  30'd    657    : data = 32'h    10871097    ;    //    auipc x1 67697      ====        auipc ra, 67697
                                                  30'd    658    : data = 32'h    01A30E33    ;    //    add x28 x6 x26      ====        add t3, t1, s10
                                                  30'd    659    : data = 32'h    009F8633    ;    //    add x12 x31 x9      ====        add a2, t6, s1
                                                  30'd    660    : data = 32'h    73298FB7    ;    //    lui x31 471704      ====        lui t6, 471704
                                                  30'd    661    : data = 32'h    09C48F93    ;    //    addi x31 x9 156      ====        addi t6, s1, 156
                                                  30'd    662    : data = 32'h    6FFE0897    ;    //    auipc x17 458720      ====        auipc a7, 458720
                                                  30'd    663    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    664    : data = 32'h    4890A0EF    ;    //    jal x1 44168      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_25
                                                  30'd    665    : data = 32'h    800008B7    ;    //    lui x17 524288      ====        li a7, 0x80000000 #start riscv_int_numeric_corner_stream_3
                                                  30'd    666    : data = 32'h    00088893    ;    //    addi x17 x17 0      ====        li a7, 0x80000000 #start riscv_int_numeric_corner_stream_3
                                                  30'd    667    : data = 32'h    FFF00B13    ;    //    addi x22 x0 -1      ====        li s6, 0xffffffff
                                                  30'd    668    : data = 32'h    80000CB7    ;    //    lui x25 524288      ====        li s9, 0x80000000
                                                  30'd    669    : data = 32'h    000C8C93    ;    //    addi x25 x25 0      ====        li s9, 0x80000000
                                                  30'd    670    : data = 32'h    FFF00613    ;    //    addi x12 x0 -1      ====        li a2, 0xffffffff
                                                  30'd    671    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff
                                                  30'd    672    : data = 32'h    FFF00813    ;    //    addi x16 x0 -1      ====        li a6, 0xffffffff
                                                  30'd    673    : data = 32'h    FFF00313    ;    //    addi x6 x0 -1      ====        li t1, 0xffffffff
                                                  30'd    674    : data = 32'h    00000493    ;    //    addi x9 x0 0      ====        li s1, 0x0
                                                  30'd    675    : data = 32'h    00000693    ;    //    addi x13 x0 0      ====        li a3, 0x0
                                                  30'd    676    : data = 32'h    FFF00B93    ;    //    addi x23 x0 -1      ====        li s7, 0xffffffff
                                                  30'd    677    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    678    : data = 32'h    D755DB97    ;    //    auipc x23 882013      ====        auipc s7, 882013
                                                  30'd    679    : data = 32'h    5C8CE337    ;    //    lui x6 379086      ====        lui t1, 379086
                                                  30'd    680    : data = 32'h    97DB8813    ;    //    addi x16 x23 -1667      ====        addi a6, s7, -1667
                                                  30'd    681    : data = 32'h    0C425497    ;    //    auipc x9 50213      ====        auipc s1, 50213
                                                  30'd    682    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    683    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    684    : data = 32'h    B55CE617    ;    //    auipc x12 742862      ====        auipc a2, 742862
                                                  30'd    685    : data = 32'h    C728F837    ;    //    lui x16 815759      ====        lui a6, 815759
                                                  30'd    686    : data = 32'h    00130CB3    ;    //    add x25 x6 x1      ====        add s9, t1, ra
                                                  30'd    687    : data = 32'h    B770CB97    ;    //    auipc x23 751372      ====        auipc s7, 751372
                                                  30'd    688    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    689    : data = 32'h    00D68BB3    ;    //    add x23 x13 x13      ====        add s7, a3, a3
                                                  30'd    690    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    691    : data = 32'h    7526CB97    ;    //    auipc x23 479852      ====        auipc s7, 479852
                                                  30'd    692    : data = 32'h    016B8CB3    ;    //    add x25 x23 x22      ====        add s9, s7, s6
                                                  30'd    693    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    694    : data = 32'h    410B8B33    ;    //    sub x22 x23 x16      ====        sub s6, s7, a6
                                                  30'd    695    : data = 32'h    1460C0B7    ;    //    lui x1 83468      ====        lui ra, 83468
                                                  30'd    696    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    697    : data = 32'h    40180833    ;    //    sub x16 x16 x1      ====        sub a6, a6, ra
                                                  30'd    698    : data = 32'h    CB9E76B7    ;    //    lui x13 834023      ====        lui a3, 834023
                                                  30'd    699    : data = 32'h    0CB34697    ;    //    auipc x13 52020      ====        auipc a3, 52020
                                                  30'd    700    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    701    : data = 32'h    0AB51B37    ;    //    lui x22 43857      ====        lui s6, 43857
                                                  30'd    702    : data = 32'h    411800B3    ;    //    sub x1 x16 x17      ====        sub ra, a6, a7
                                                  30'd    703    : data = 32'h    410808B3    ;    //    sub x17 x16 x16      ====        sub a7, a6, a6
                                                  30'd    704    : data = 32'h    00C80B33    ;    //    add x22 x16 x12      ====        add s6, a6, a2
                                                  30'd    705    : data = 32'h    3E50A0EF    ;    //    jal x1 44004      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_3
                                                  30'd    706    : data = 32'h    FFF00C13    ;    //    addi x24 x0 -1      ====        li s8, 0xffffffff #start riscv_int_numeric_corner_stream_35
                                                  30'd    707    : data = 32'h    00000693    ;    //    addi x13 x0 0      ====        li a3, 0x0
                                                  30'd    708    : data = 32'h    80000437    ;    //    lui x8 524288      ====        li s0, 0x80000000
                                                  30'd    709    : data = 32'h    00040413    ;    //    addi x8 x8 0      ====        li s0, 0x80000000
                                                  30'd    710    : data = 32'h    FFF00113    ;    //    addi x2 x0 -1      ====        li sp, 0xffffffff
                                                  30'd    711    : data = 32'h    00000993    ;    //    addi x19 x0 0      ====        li s3, 0x0
                                                  30'd    712    : data = 32'h    FFF00913    ;    //    addi x18 x0 -1      ====        li s2, 0xffffffff
                                                  30'd    713    : data = 32'h    83C533B7    ;    //    lui x7 539731      ====        li t2, 0x83c5299f
                                                  30'd    714    : data = 32'h    99F38393    ;    //    addi x7 x7 -1633      ====        li t2, 0x83c5299f
                                                  30'd    715    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff
                                                  30'd    716    : data = 32'h    FFF00493    ;    //    addi x9 x0 -1      ====        li s1, 0xffffffff
                                                  30'd    717    : data = 32'h    00000E13    ;    //    addi x28 x0 0      ====        li t3, 0x0
                                                  30'd    718    : data = 32'h    05FE0413    ;    //    addi x8 x28 95      ====        addi s0, t3, 95
                                                  30'd    719    : data = 32'h    40D98E33    ;    //    sub x28 x19 x13      ====        sub t3, s3, a3
                                                  30'd    720    : data = 32'h    ED364497    ;    //    auipc x9 971620      ====        auipc s1, 971620
                                                  30'd    721    : data = 32'h    B65B2417    ;    //    auipc x8 746930      ====        auipc s0, 746930
                                                  30'd    722    : data = 32'h    FA763C37    ;    //    lui x24 1025891      ====        lui s8, 1025891
                                                  30'd    723    : data = 32'h    41CE0433    ;    //    sub x8 x28 x28      ====        sub s0, t3, t3
                                                  30'd    724    : data = 32'h    402980B3    ;    //    sub x1 x19 x2      ====        sub ra, s3, sp
                                                  30'd    725    : data = 32'h    02E98693    ;    //    addi x13 x19 46      ====        addi a3, s3, 46
                                                  30'd    726    : data = 32'h    93FD2E37    ;    //    lui x28 606162      ====        lui t3, 606162
                                                  30'd    727    : data = 32'h    0B046137    ;    //    lui x2 45126      ====        lui sp, 45126
                                                  30'd    728    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    729    : data = 32'h    013983B3    ;    //    add x7 x19 x19      ====        add t2, s3, s3
                                                  30'd    730    : data = 32'h    41238C33    ;    //    sub x24 x7 x18      ====        sub s8, t2, s2
                                                  30'd    731    : data = 32'h    1C319137    ;    //    lui x2 115481      ====        lui sp, 115481
                                                  30'd    732    : data = 32'h    41238E33    ;    //    sub x28 x7 x18      ====        sub t3, t2, s2
                                                  30'd    733    : data = 32'h    A9208993    ;    //    addi x19 x1 -1390      ====        addi s3, ra, -1390
                                                  30'd    734    : data = 32'h    01CC09B3    ;    //    add x19 x24 x28      ====        add s3, s8, t3
                                                  30'd    735    : data = 32'h    1CD19E37    ;    //    lui x28 118041      ====        lui t3, 118041
                                                  30'd    736    : data = 32'h    3FC38913    ;    //    addi x18 x7 1020      ====        addi s2, t2, 1020
                                                  30'd    737    : data = 32'h    780F7E37    ;    //    lui x28 491767      ====        lui t3, 491767
                                                  30'd    738    : data = 32'h    E0298693    ;    //    addi x13 x19 -510      ====        addi a3, s3, -510
                                                  30'd    739    : data = 32'h    40248133    ;    //    sub x2 x9 x2      ====        sub sp, s1, sp
                                                  30'd    740    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    741    : data = 32'h    007983B3    ;    //    add x7 x19 x7      ====        add t2, s3, t2
                                                  30'd    742    : data = 32'h    947F1E37    ;    //    lui x28 608241      ====        lui t3, 608241
                                                  30'd    743    : data = 32'h    01290433    ;    //    add x8 x18 x18      ====        add s0, s2, s2
                                                  30'd    744    : data = 32'h    C106AE37    ;    //    lui x28 790634      ====        lui t3, 790634
                                                  30'd    745    : data = 32'h    3450A0EF    ;    //    jal x1 43844      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_35
                                                  30'd    746    : data = 32'h    00B4C7B7    ;    //    lui x15 2892      ====        li a5, 0xb4c19b #start riscv_int_numeric_corner_stream_15
                                                  30'd    747    : data = 32'h    19B78793    ;    //    addi x15 x15 411      ====        li a5, 0xb4c19b #start riscv_int_numeric_corner_stream_15
                                                  30'd    748    : data = 32'h    80000437    ;    //    lui x8 524288      ====        li s0, 0x80000000
                                                  30'd    749    : data = 32'h    00040413    ;    //    addi x8 x8 0      ====        li s0, 0x80000000
                                                  30'd    750    : data = 32'h    00000E13    ;    //    addi x28 x0 0      ====        li t3, 0x0
                                                  30'd    751    : data = 32'h    80000737    ;    //    lui x14 524288      ====        li a4, 0x80000000
                                                  30'd    752    : data = 32'h    00070713    ;    //    addi x14 x14 0      ====        li a4, 0x80000000
                                                  30'd    753    : data = 32'h    00000093    ;    //    addi x1 x0 0      ====        li ra, 0x0
                                                  30'd    754    : data = 32'h    FFF00693    ;    //    addi x13 x0 -1      ====        li a3, 0xffffffff
                                                  30'd    755    : data = 32'h    FFF00893    ;    //    addi x17 x0 -1      ====        li a7, 0xffffffff
                                                  30'd    756    : data = 32'h    96D13AB7    ;    //    lui x21 617747      ====        li s5, 0x96d12823
                                                  30'd    757    : data = 32'h    823A8A93    ;    //    addi x21 x21 -2013      ====        li s5, 0x96d12823
                                                  30'd    758    : data = 32'h    80000CB7    ;    //    lui x25 524288      ====        li s9, 0x80000000
                                                  30'd    759    : data = 32'h    000C8C93    ;    //    addi x25 x25 0      ====        li s9, 0x80000000
                                                  30'd    760    : data = 32'h    800003B7    ;    //    lui x7 524288      ====        li t2, 0x80000000
                                                  30'd    761    : data = 32'h    00038393    ;    //    addi x7 x7 0      ====        li t2, 0x80000000
                                                  30'd    762    : data = 32'h    40F083B3    ;    //    sub x7 x1 x15      ====        sub t2, ra, a5
                                                  30'd    763    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    764    : data = 32'h    001C87B3    ;    //    add x15 x25 x1      ====        add a5, s9, ra
                                                  30'd    765    : data = 32'h    A53CB797    ;    //    auipc x15 676811      ====        auipc a5, 676811
                                                  30'd    766    : data = 32'h    58ADE437    ;    //    lui x8 363230      ====        lui s0, 363230
                                                  30'd    767    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    768    : data = 32'h    F5039AB7    ;    //    lui x21 1003577      ====        lui s5, 1003577
                                                  30'd    769    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    770    : data = 32'h    C1EC8E13    ;    //    addi x28 x25 -994      ====        addi t3, s9, -994
                                                  30'd    771    : data = 32'h    2C7716B7    ;    //    lui x13 182129      ====        lui a3, 182129
                                                  30'd    772    : data = 32'h    9F0D3C97    ;    //    auipc x25 651475      ====        auipc s9, 651475
                                                  30'd    773    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    774    : data = 32'h    00FA8733    ;    //    add x14 x21 x15      ====        add a4, s5, a5
                                                  30'd    775    : data = 32'h    A1438713    ;    //    addi x14 x7 -1516      ====        addi a4, t2, -1516
                                                  30'd    776    : data = 32'h    367F0797    ;    //    auipc x15 223216      ====        auipc a5, 223216
                                                  30'd    777    : data = 32'h    00D08733    ;    //    add x14 x1 x13      ====        add a4, ra, a3
                                                  30'd    778    : data = 32'h    5F0CCCB7    ;    //    lui x25 389324      ====        lui s9, 389324
                                                  30'd    779    : data = 32'h    F25343B7    ;    //    lui x7 992564      ====        lui t2, 992564
                                                  30'd    780    : data = 32'h    00F086B3    ;    //    add x13 x1 x15      ====        add a3, ra, a5
                                                  30'd    781    : data = 32'h    B7212437    ;    //    lui x8 750098      ====        lui s0, 750098
                                                  30'd    782    : data = 32'h    2B10A0EF    ;    //    jal x1 43696      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_15
                                                  30'd    783    : data = 32'h    80000937    ;    //    lui x18 524288      ====        li s2, 0x80000000 #start riscv_int_numeric_corner_stream_13
                                                  30'd    784    : data = 32'h    00090913    ;    //    addi x18 x18 0      ====        li s2, 0x80000000 #start riscv_int_numeric_corner_stream_13
                                                  30'd    785    : data = 32'h    800008B7    ;    //    lui x17 524288      ====        li a7, 0x80000000
                                                  30'd    786    : data = 32'h    00088893    ;    //    addi x17 x17 0      ====        li a7, 0x80000000
                                                  30'd    787    : data = 32'h    80000CB7    ;    //    lui x25 524288      ====        li s9, 0x80000000
                                                  30'd    788    : data = 32'h    000C8C93    ;    //    addi x25 x25 0      ====        li s9, 0x80000000
                                                  30'd    789    : data = 32'h    00000C13    ;    //    addi x24 x0 0      ====        li s8, 0x0
                                                  30'd    790    : data = 32'h    00000313    ;    //    addi x6 x0 0      ====        li t1, 0x0
                                                  30'd    791    : data = 32'h    DC5AFDB7    ;    //    lui x27 902575      ====        li s11, 0xdc5af53e
                                                  30'd    792    : data = 32'h    53ED8D93    ;    //    addi x27 x27 1342      ====        li s11, 0xdc5af53e
                                                  30'd    793    : data = 32'h    00000793    ;    //    addi x15 x0 0      ====        li a5, 0x0
                                                  30'd    794    : data = 32'h    FFF00093    ;    //    addi x1 x0 -1      ====        li ra, 0xffffffff
                                                  30'd    795    : data = 32'h    00000F93    ;    //    addi x31 x0 0      ====        li t6, 0x0
                                                  30'd    796    : data = 32'h    6DDF0A37    ;    //    lui x20 450032      ====        li s4, 0x6ddefb74
                                                  30'd    797    : data = 32'h    B74A0A13    ;    //    addi x20 x20 -1164      ====        li s4, 0x6ddefb74
                                                  30'd    798    : data = 32'h    41BC0A33    ;    //    sub x20 x24 x27      ====        sub s4, s8, s11
                                                  30'd    799    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    800    : data = 32'h    411C07B3    ;    //    sub x15 x24 x17      ====        sub a5, s8, a7
                                                  30'd    801    : data = 32'h    01B880B3    ;    //    add x1 x17 x27      ====        add ra, a7, s11
                                                  30'd    802    : data = 32'h    E8A57C17    ;    //    auipc x24 952919      ====        auipc s8, 952919
                                                  30'd    803    : data = 32'h    5ADD3C97    ;    //    auipc x25 372179      ====        auipc s9, 372179
                                                  30'd    804    : data = 32'h    7B55C337    ;    //    lui x6 505180      ====        lui t1, 505180
                                                  30'd    805    : data = 32'h    01BD8C33    ;    //    add x24 x27 x27      ====        add s8, s11, s11
                                                  30'd    806    : data = 32'h    931D2C17    ;    //    auipc x24 602578      ====        auipc s8, 602578
                                                  30'd    807    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    808    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    809    : data = 32'h    24434317    ;    //    auipc x6 148532      ====        auipc t1, 148532
                                                  30'd    810    : data = 32'h    AD350DB7    ;    //    lui x27 709456      ====        lui s11, 709456
                                                  30'd    811    : data = 32'h    A72C8C93    ;    //    addi x25 x25 -1422      ====        addi s9, s9, -1422
                                                  30'd    812    : data = 32'h    67CD8913    ;    //    addi x18 x27 1660      ====        addi s2, s11, 1660
                                                  30'd    813    : data = 32'h    01878CB3    ;    //    add x25 x15 x24      ====        add s9, a5, s8
                                                  30'd    814    : data = 32'h    CBC78797    ;    //    auipc x15 834680      ====        auipc a5, 834680
                                                  30'd    815    : data = 32'h    018880B3    ;    //    add x1 x17 x24      ====        add ra, a7, s8
                                                  30'd    816    : data = 32'h    B6BA2CB7    ;    //    lui x25 748450      ====        lui s9, 748450
                                                  30'd    817    : data = 32'h    41990CB3    ;    //    sub x25 x18 x25      ====        sub s9, s2, s9
                                                  30'd    818    : data = 32'h    D71C0313    ;    //    addi x6 x24 -655      ====        addi t1, s8, -655
                                                  30'd    819    : data = 32'h    CC130D93    ;    //    addi x27 x6 -831      ====        addi s11, t1, -831
                                                  30'd    820    : data = 32'h    6E9B9F97    ;    //    auipc x31 453049      ====        auipc t6, 453049
                                                  30'd    821    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    822    : data = 32'h    0AB5ADB7    ;    //    lui x27 43866      ====        lui s11, 43866
                                                  30'd    823    : data = 32'h    D6CD8A13    ;    //    addi x20 x27 -660      ====        addi s4, s11, -660
                                                  30'd    824    : data = 32'h    40F78A33    ;    //    sub x20 x15 x15      ====        sub s4, a5, a5
                                                  30'd    825    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    826    : data = 32'h    DD4B8A37    ;    //    lui x20 906424      ====        lui s4, 906424
                                                  30'd    827    : data = 32'h    1FD0A0EF    ;    //    jal x1 43516      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_13
                                                  30'd    828    : data = 32'h    0EF34CB7    ;    //    lui x25 61236      ====        li s9, 0xef34712 #start riscv_int_numeric_corner_stream_33
                                                  30'd    829    : data = 32'h    712C8C93    ;    //    addi x25 x25 1810      ====        li s9, 0xef34712 #start riscv_int_numeric_corner_stream_33
                                                  30'd    830    : data = 32'h    800002B7    ;    //    lui x5 524288      ====        li t0, 0x80000000
                                                  30'd    831    : data = 32'h    00028293    ;    //    addi x5 x5 0      ====        li t0, 0x80000000
                                                  30'd    832    : data = 32'h    00000493    ;    //    addi x9 x0 0      ====        li s1, 0x0
                                                  30'd    833    : data = 32'h    FFF00D93    ;    //    addi x27 x0 -1      ====        li s11, 0xffffffff
                                                  30'd    834    : data = 32'h    FFF00813    ;    //    addi x16 x0 -1      ====        li a6, 0xffffffff
                                                  30'd    835    : data = 32'h    FFF00913    ;    //    addi x18 x0 -1      ====        li s2, 0xffffffff
                                                  30'd    836    : data = 32'h    00000E93    ;    //    addi x29 x0 0      ====        li t4, 0x0
                                                  30'd    837    : data = 32'h    FFF00B93    ;    //    addi x23 x0 -1      ====        li s7, 0xffffffff
                                                  30'd    838    : data = 32'h    FFF00D13    ;    //    addi x26 x0 -1      ====        li s10, 0xffffffff
                                                  30'd    839    : data = 32'h    FFF00413    ;    //    addi x8 x0 -1      ====        li s0, 0xffffffff
                                                  30'd    840    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    841    : data = 32'h    D8DDFD97    ;    //    auipc x27 888287      ====        auipc s11, 888287
                                                  30'd    842    : data = 32'h    F9490293    ;    //    addi x5 x18 -108      ====        addi t0, s2, -108
                                                  30'd    843    : data = 32'h    01D48433    ;    //    add x8 x9 x29      ====        add s0, s1, t4
                                                  30'd    844    : data = 32'h    1C7D8913    ;    //    addi x18 x27 455      ====        addi s2, s11, 455
                                                  30'd    845    : data = 32'h    95248D93    ;    //    addi x27 x9 -1710      ====        addi s11, s1, -1710
                                                  30'd    846    : data = 32'h    41A40CB3    ;    //    sub x25 x8 x26      ====        sub s9, s0, s10
                                                  30'd    847    : data = 32'h    409E8933    ;    //    sub x18 x29 x9      ====        sub s2, t4, s1
                                                  30'd    848    : data = 32'h    95EB8813    ;    //    addi x16 x23 -1698      ====        addi a6, s7, -1698
                                                  30'd    849    : data = 32'h    00540DB3    ;    //    add x27 x8 x5      ====        add s11, s0, t0
                                                  30'd    850    : data = 32'h    FBAB8D93    ;    //    addi x27 x23 -70      ====        addi s11, s7, -70
                                                  30'd    851    : data = 32'h    1D848B93    ;    //    addi x23 x9 472      ====        addi s7, s1, 472
                                                  30'd    852    : data = 32'h    46A90493    ;    //    addi x9 x18 1130      ====        addi s1, s2, 1130
                                                  30'd    853    : data = 32'h    DBFD8913    ;    //    addi x18 x27 -577      ====        addi s2, s11, -577
                                                  30'd    854    : data = 32'h    00828BB3    ;    //    add x23 x5 x8      ====        add s7, t0, s0
                                                  30'd    855    : data = 32'h    BD3D6417    ;    //    auipc x8 775126      ====        auipc s0, 775126
                                                  30'd    856    : data = 32'h    412D0BB3    ;    //    sub x23 x26 x18      ====        sub s7, s10, s2
                                                  30'd    857    : data = 32'h    DBB8A817    ;    //    auipc x16 899978      ====        auipc a6, 899978
                                                  30'd    858    : data = 32'h    9C1B8493    ;    //    addi x9 x23 -1599      ====        addi s1, s7, -1599
                                                  30'd    859    : data = 32'h    E2290413    ;    //    addi x8 x18 -478      ====        addi s0, s2, -478
                                                  30'd    860    : data = 32'h    01BE8D33    ;    //    add x26 x29 x27      ====        add s10, t4, s11
                                                  30'd    861    : data = 32'h    218F1CB7    ;    //    lui x25 137457      ====        lui s9, 137457
                                                  30'd    862    : data = 32'h    1710A0EF    ;    //    jal x1 43376      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_33
                                                  30'd    863    : data = 32'h    0AFAA1B7    ;    //    lui x3 44970      ====        li gp, 0xafaa20e #start riscv_int_numeric_corner_stream_36
                                                  30'd    864    : data = 32'h    20E18193    ;    //    addi x3 x3 526      ====        li gp, 0xafaa20e #start riscv_int_numeric_corner_stream_36
                                                  30'd    865    : data = 32'h    7B54B7B7    ;    //    lui x15 505163      ====        li a5, 0x7b54b34b
                                                  30'd    866    : data = 32'h    34B78793    ;    //    addi x15 x15 843      ====        li a5, 0x7b54b34b
                                                  30'd    867    : data = 32'h    13152BB7    ;    //    lui x23 78162      ====        li s7, 0x13152550
                                                  30'd    868    : data = 32'h    550B8B93    ;    //    addi x23 x23 1360      ====        li s7, 0x13152550
                                                  30'd    869    : data = 32'h    00000813    ;    //    addi x16 x0 0      ====        li a6, 0x0
                                                  30'd    870    : data = 32'h    80000B37    ;    //    lui x22 524288      ====        li s6, 0x80000000
                                                  30'd    871    : data = 32'h    000B0B13    ;    //    addi x22 x22 0      ====        li s6, 0x80000000
                                                  30'd    872    : data = 32'h    00000313    ;    //    addi x6 x0 0      ====        li t1, 0x0
                                                  30'd    873    : data = 32'h    FFF00C13    ;    //    addi x24 x0 -1      ====        li s8, 0xffffffff
                                                  30'd    874    : data = 32'h    00000C93    ;    //    addi x25 x0 0      ====        li s9, 0x0
                                                  30'd    875    : data = 32'h    00000993    ;    //    addi x19 x0 0      ====        li s3, 0x0
                                                  30'd    876    : data = 32'h    FFF00613    ;    //    addi x12 x0 -1      ====        li a2, 0xffffffff
                                                  30'd    877    : data = 32'h    017307B3    ;    //    add x15 x6 x23      ====        add a5, t1, s7
                                                  30'd    878    : data = 32'h    00F98B33    ;    //    add x22 x19 x15      ====        add s6, s3, a5
                                                  30'd    879    : data = 32'h    1C746B97    ;    //    auipc x23 116550      ====        auipc s7, 116550
                                                  30'd    880    : data = 32'h    00FC8BB3    ;    //    add x23 x25 x15      ====        add s7, s9, a5
                                                  30'd    881    : data = 32'h    CA3401B7    ;    //    lui x3 828224      ====        lui gp, 828224
                                                  30'd    882    : data = 32'h    418C07B3    ;    //    sub x15 x24 x24      ====        sub a5, s8, s8
                                                  30'd    883    : data = 32'h    41678833    ;    //    sub x16 x15 x22      ====        sub a6, a5, s6
                                                  30'd    884    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    885    : data = 32'h    003C87B3    ;    //    add x15 x25 x3      ====        add a5, s9, gp
                                                  30'd    886    : data = 32'h    403B0BB3    ;    //    sub x23 x22 x3      ====        sub s7, s6, gp
                                                  30'd    887    : data = 32'h    010C8CB3    ;    //    add x25 x25 x16      ====        add s9, s9, a6
                                                  30'd    888    : data = 32'h    01030833    ;    //    add x16 x6 x16      ====        add a6, t1, a6
                                                  30'd    889    : data = 32'h    41618C33    ;    //    sub x24 x3 x22      ====        sub s8, gp, s6
                                                  30'd    890    : data = 32'h    03333C37    ;    //    lui x24 13107      ====        lui s8, 13107
                                                  30'd    891    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    892    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    893    : data = 32'h    41618CB3    ;    //    sub x25 x3 x22      ====        sub s9, gp, s6
                                                  30'd    894    : data = 32'h    41730833    ;    //    sub x16 x6 x23      ====        sub a6, t1, s7
                                                  30'd    895    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    896    : data = 32'h    585B4637    ;    //    lui x12 361908      ====        lui a2, 361908
                                                  30'd    897    : data = 32'h    00378CB3    ;    //    add x25 x15 x3      ====        add s9, a5, gp
                                                  30'd    898    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    899    : data = 32'h    512C0C93    ;    //    addi x25 x24 1298      ====        addi s9, s8, 1298
                                                  30'd    900    : data = 32'h    87AA5997    ;    //    auipc x19 555685      ====        auipc s3, 555685
                                                  30'd    901    : data = 32'h    418C0BB3    ;    //    sub x23 x24 x24      ====        sub s7, s8, s8
                                                  30'd    902    : data = 32'h    016B0CB3    ;    //    add x25 x22 x22      ====        add s9, s6, s6
                                                  30'd    903    : data = 32'h    013B0333    ;    //    add x6 x22 x19      ====        add t1, s6, s3
                                                  30'd    904    : data = 32'h    0C90A0EF    ;    //    jal x1 43208      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_36
                                                  30'd    905    : data = 32'h    80000937    ;    //    lui x18 524288      ====        li s2, 0x80000000 #start riscv_int_numeric_corner_stream_19
                                                  30'd    906    : data = 32'h    00090913    ;    //    addi x18 x18 0      ====        li s2, 0x80000000 #start riscv_int_numeric_corner_stream_19
                                                  30'd    907    : data = 32'h    5FA92837    ;    //    lui x16 391826      ====        li a6, 0x5fa92591
                                                  30'd    908    : data = 32'h    59180813    ;    //    addi x16 x16 1425      ====        li a6, 0x5fa92591
                                                  30'd    909    : data = 32'h    00000893    ;    //    addi x17 x0 0      ====        li a7, 0x0
                                                  30'd    910    : data = 32'h    00000693    ;    //    addi x13 x0 0      ====        li a3, 0x0
                                                  30'd    911    : data = 32'h    EE38F0B7    ;    //    lui x1 975759      ====        li ra, 0xee38ef7f
                                                  30'd    912    : data = 32'h    F7F08093    ;    //    addi x1 x1 -129      ====        li ra, 0xee38ef7f
                                                  30'd    913    : data = 32'h    80000DB7    ;    //    lui x27 524288      ====        li s11, 0x80000000
                                                  30'd    914    : data = 32'h    000D8D93    ;    //    addi x27 x27 0      ====        li s11, 0x80000000
                                                  30'd    915    : data = 32'h    FFF00493    ;    //    addi x9 x0 -1      ====        li s1, 0xffffffff
                                                  30'd    916    : data = 32'h    80000E37    ;    //    lui x28 524288      ====        li t3, 0x80000000
                                                  30'd    917    : data = 32'h    000E0E13    ;    //    addi x28 x28 0      ====        li t3, 0x80000000
                                                  30'd    918    : data = 32'h    80000137    ;    //    lui x2 524288      ====        li sp, 0x80000000
                                                  30'd    919    : data = 32'h    00010113    ;    //    addi x2 x2 0      ====        li sp, 0x80000000
                                                  30'd    920    : data = 32'h    00000D13    ;    //    addi x26 x0 0      ====        li s10, 0x0
                                                  30'd    921    : data = 32'h    59490093    ;    //    addi x1 x18 1428      ====        addi ra, s2, 1428
                                                  30'd    922    : data = 32'h    412D0E33    ;    //    sub x28 x26 x18      ====        sub t3, s10, s2
                                                  30'd    923    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    924    : data = 32'h    41B800B3    ;    //    sub x1 x16 x27      ====        sub ra, a6, s11
                                                  30'd    925    : data = 32'h    01208933    ;    //    add x18 x1 x18      ====        add s2, ra, s2
                                                  30'd    926    : data = 32'h    F9986DB7    ;    //    lui x27 1022342      ====        lui s11, 1022342
                                                  30'd    927    : data = 32'h    B44FE117    ;    //    auipc x2 738558      ====        auipc sp, 738558
                                                  30'd    928    : data = 32'h    958AD0B7    ;    //    lui x1 612525      ====        lui ra, 612525
                                                  30'd    929    : data = 32'h    2A197E17    ;    //    auipc x28 172439      ====        auipc t3, 172439
                                                  30'd    930    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    931    : data = 32'h    36908E13    ;    //    addi x28 x1 873      ====        addi t3, ra, 873
                                                  30'd    932    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    933    : data = 32'h    F7E0E0B7    ;    //    lui x1 1015310      ====        lui ra, 1015310
                                                  30'd    934    : data = 32'h    604816B7    ;    //    lui x13 394369      ====        lui a3, 394369
                                                  30'd    935    : data = 32'h    012D80B3    ;    //    add x1 x27 x18      ====        add ra, s11, s2
                                                  30'd    936    : data = 32'h    ABFD0813    ;    //    addi x16 x26 -1345      ====        addi a6, s10, -1345
                                                  30'd    937    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    938    : data = 32'h    58B3FD97    ;    //    auipc x27 363327      ====        auipc s11, 363327
                                                  30'd    939    : data = 32'h    00908DB3    ;    //    add x27 x1 x9      ====        add s11, ra, s1
                                                  30'd    940    : data = 32'h    83643E17    ;    //    auipc x28 538179      ====        auipc t3, 538179
                                                  30'd    941    : data = 32'h    0350A0EF    ;    //    jal x1 43060      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_19
                                                  30'd    942    : data = 32'h    FFF00D93    ;    //    addi x27 x0 -1      ====        li s11, 0xffffffff #start riscv_int_numeric_corner_stream_2
                                                  30'd    943    : data = 32'h    213EC5B7    ;    //    lui x11 136172      ====        li a1, 0x213ec4a9
                                                  30'd    944    : data = 32'h    4A958593    ;    //    addi x11 x11 1193      ====        li a1, 0x213ec4a9
                                                  30'd    945    : data = 32'h    00000293    ;    //    addi x5 x0 0      ====        li t0, 0x0
                                                  30'd    946    : data = 32'h    00000613    ;    //    addi x12 x0 0      ====        li a2, 0x0
                                                  30'd    947    : data = 32'h    C1F611B7    ;    //    lui x3 794465      ====        li gp, 0xc1f61669
                                                  30'd    948    : data = 32'h    66918193    ;    //    addi x3 x3 1641      ====        li gp, 0xc1f61669
                                                  30'd    949    : data = 32'h    FFF00393    ;    //    addi x7 x0 -1      ====        li t2, 0xffffffff
                                                  30'd    950    : data = 32'h    80000137    ;    //    lui x2 524288      ====        li sp, 0x80000000
                                                  30'd    951    : data = 32'h    00010113    ;    //    addi x2 x2 0      ====        li sp, 0x80000000
                                                  30'd    952    : data = 32'h    80000AB7    ;    //    lui x21 524288      ====        li s5, 0x80000000
                                                  30'd    953    : data = 32'h    000A8A93    ;    //    addi x21 x21 0      ====        li s5, 0x80000000
                                                  30'd    954    : data = 32'h    800007B7    ;    //    lui x15 524288      ====        li a5, 0x80000000
                                                  30'd    955    : data = 32'h    00078793    ;    //    addi x15 x15 0      ====        li a5, 0x80000000
                                                  30'd    956    : data = 32'h    00000E13    ;    //    addi x28 x0 0      ====        li t3, 0x0
                                                  30'd    957    : data = 32'h    4C1C1A97    ;    //    auipc x21 311745      ====        auipc s5, 311745
                                                  30'd    958    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    959    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    960    : data = 32'h    CA378E13    ;    //    addi x28 x15 -861      ====        addi t3, a5, -861
                                                  30'd    961    : data = 32'h    41B107B3    ;    //    sub x15 x2 x27      ====        sub a5, sp, s11
                                                  30'd    962    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    963    : data = 32'h    6CCE9E37    ;    //    lui x28 445673      ====        lui t3, 445673
                                                  30'd    964    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    965    : data = 32'h    C0F02DB7    ;    //    lui x27 790274      ====        lui s11, 790274
                                                  30'd    966    : data = 32'h    40C60DB3    ;    //    sub x27 x12 x12      ====        sub s11, a2, a2
                                                  30'd    967    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    968    : data = 32'h    402E02B3    ;    //    sub x5 x28 x2      ====        sub t0, t3, sp
                                                  30'd    969    : data = 32'h    1C13AE17    ;    //    auipc x28 115002      ====        auipc t3, 115002
                                                  30'd    970    : data = 32'h    D92D6197    ;    //    auipc x3 889558      ====        auipc gp, 889558
                                                  30'd    971    : data = 32'h    FF50C637    ;    //    lui x12 1045772      ====        lui a2, 1045772
                                                  30'd    972    : data = 32'h    003A81B3    ;    //    add x3 x21 x3      ====        add gp, s5, gp
                                                  30'd    973    : data = 32'h    864A07B7    ;    //    lui x15 550048      ====        lui a5, 550048
                                                  30'd    974    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    975    : data = 32'h    EF9145B7    ;    //    lui x11 981268      ====        lui a1, 981268
                                                  30'd    976    : data = 32'h    00FE2E37    ;    //    lui x28 4066      ====        lui t3, 4066
                                                  30'd    977    : data = 32'h    EB118E13    ;    //    addi x28 x3 -335      ====        addi t3, gp, -335
                                                  30'd    978    : data = 32'h    015787B3    ;    //    add x15 x15 x21      ====        add a5, a5, s5
                                                  30'd    979    : data = 32'h    F824A137    ;    //    lui x2 1016394      ====        lui sp, 1016394
                                                  30'd    980    : data = 32'h    7980A0EF    ;    //    jal x1 42904      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_2
                                                  30'd    981    : data = 32'h    019DD713    ;    //    srli x14 x27 25      ====        srli a4, s11, 25
                                                  30'd    982    : data = 32'h    018CCC33    ;    //    xor x24 x25 x24      ====        xor s8, s9, s8
                                                  30'd    983    : data = 32'h    BCA66713    ;    //    ori x14 x12 -1078      ====        ori a4, a2, -1078
                                                  30'd    984    : data = 32'h    00AAF3B3    ;    //    and x7 x21 x10      ====        and t2, s5, a0
                                                  30'd    985    : data = 32'h    00339913    ;    //    slli x18 x7 3      ====        slli s2, t2, 3
                                                  30'd    986    : data = 32'h    412CD693    ;    //    srai x13 x25 18      ====        srai a3, s9, 18
                                                  30'd    987    : data = 32'h    006F3733    ;    //    sltu x14 x30 x6      ====        sltu a4, t5, t1
                                                  30'd    988    : data = 32'h    41B2DEB3    ;    //    sra x29 x5 x27      ====        sra t4, t0, s11
                                                  30'd    989    : data = 32'h    94F4EBB7    ;    //    lui x23 610126      ====        lui s7, 610126
                                                  30'd    990    : data = 32'h    C3AC4713    ;    //    xori x14 x24 -966      ====        xori a4, s8, -966
                                                  30'd    991    : data = 32'h    97FB0817    ;    //    auipc x16 622512      ====        auipc a6, 622512
                                                  30'd    992    : data = 32'h    CFA81197    ;    //    auipc x3 850561      ====        auipc gp, 850561
                                                  30'd    993    : data = 32'h    9C636013    ;    //    ori x0 x6 -1594      ====        ori zero, t1, -1594
                                                  30'd    994    : data = 32'h    928B2093    ;    //    slti x1 x22 -1752      ====        slti ra, s6, -1752
                                                  30'd    995    : data = 32'h    00CFFDB3    ;    //    and x27 x31 x12      ====        and s11, t6, a2
                                                  30'd    996    : data = 32'h    01881BB3    ;    //    sll x23 x16 x24      ====        sll s7, a6, s8
                                                  30'd    997    : data = 32'h    7C05ED93    ;    //    ori x27 x11 1984      ====        ori s11, a1, 1984
                                                  30'd    998    : data = 32'h    41A555B3    ;    //    sra x11 x10 x26      ====        sra a1, a0, s10
                                                  30'd    999    : data = 32'h    0435E093    ;    //    ori x1 x11 67      ====        ori ra, a1, 67
                                                  30'd    1000    : data = 32'h    01BAC0B3    ;    //    xor x1 x21 x27      ====        xor ra, s5, s11
                                                  30'd    1001    : data = 32'h    01CB58B3    ;    //    srl x17 x22 x28      ====        srl a7, s6, t3
                                                  30'd    1002    : data = 32'h    70A60B93    ;    //    addi x23 x12 1802      ====        addi s7, a2, 1802
                                                  30'd    1003    : data = 32'h    01544933    ;    //    xor x18 x8 x21      ====        xor s2, s0, s5
                                                  30'd    1004    : data = 32'h    4103DB33    ;    //    sra x22 x7 x16      ====        sra s6, t2, a6
                                                  30'd    1005    : data = 32'h    017D2DB3    ;    //    slt x27 x26 x23      ====        slt s11, s10, s7
                                                  30'd    1006    : data = 32'h    00A782B3    ;    //    add x5 x15 x10      ====        add t0, a5, a0
                                                  30'd    1007    : data = 32'h    DABFF413    ;    //    andi x8 x31 -597      ====        andi s0, t6, -597
                                                  30'd    1008    : data = 32'h    4116D913    ;    //    srai x18 x13 17      ====        srai s2, a3, 17
                                                  30'd    1009    : data = 32'h    0128E1B3    ;    //    or x3 x17 x18      ====        or gp, a7, s2
                                                  30'd    1010    : data = 32'h    01CD39B3    ;    //    sltu x19 x26 x28      ====        sltu s3, s10, t3
                                                  30'd    1011    : data = 32'h    004FD613    ;    //    srli x12 x31 4      ====        srli a2, t6, 4
                                                  30'd    1012    : data = 32'h    0053D0B3    ;    //    srl x1 x7 x5      ====        srl ra, t2, t0
                                                  30'd    1013    : data = 32'h    011E2FB3    ;    //    slt x31 x28 x17      ====        slt t6, t3, a7
                                                  30'd    1014    : data = 32'h    00C582B3    ;    //    add x5 x11 x12      ====        add t0, a1, a2
                                                  30'd    1015    : data = 32'h    88A98B97    ;    //    auipc x23 559768      ====        auipc s7, 559768
                                                  30'd    1016    : data = 32'h    01732733    ;    //    slt x14 x6 x23      ====        slt a4, t1, s7
                                                  30'd    1017    : data = 32'h    D0C34D13    ;    //    xori x26 x6 -756      ====        xori s10, t1, -756
                                                  30'd    1018    : data = 32'h    ADCEC693    ;    //    xori x13 x29 -1316      ====        xori a3, t4, -1316
                                                  30'd    1019    : data = 32'h    40DD5933    ;    //    sra x18 x26 x13      ====        sra s2, s10, a3
                                                  30'd    1020    : data = 32'h    8B1F6317    ;    //    auipc x6 569846      ====        auipc t1, 569846
                                                  30'd    1021    : data = 32'h    00C2A833    ;    //    slt x16 x5 x12      ====        slt a6, t0, a2
                                                  30'd    1022    : data = 32'h    00425033    ;    //    srl x0 x4 x4      ====        srl zero, tp, tp
                                                  30'd    1023    : data = 32'h    003E06B3    ;    //    add x13 x28 x3      ====        add a3, t3, gp
                                                  30'd    1024    : data = 32'h    01E617B3    ;    //    sll x15 x12 x30      ====        sll a5, a2, t5
                                                  30'd    1025    : data = 32'h    010F30B3    ;    //    sltu x1 x30 x16      ====        sltu ra, t5, a6
                                                  30'd    1026    : data = 32'h    B0E0E837    ;    //    lui x16 724494      ====        lui a6, 724494
                                                  30'd    1027    : data = 32'h    F6972E13    ;    //    slti x28 x14 -151      ====        slti t3, a4, -151
                                                  30'd    1028    : data = 32'h    A00E2793    ;    //    slti x15 x28 -1536      ====        slti a5, t3, -1536
                                                  30'd    1029    : data = 32'h    C2E47493    ;    //    andi x9 x8 -978      ====        andi s1, s0, -978
                                                  30'd    1030    : data = 32'h    5956D437    ;    //    lui x8 365933      ====        lui s0, 365933
                                                  30'd    1031    : data = 32'h    00BDE733    ;    //    or x14 x27 x11      ====        or a4, s11, a1
                                                  30'd    1032    : data = 32'h    E8C2F937    ;    //    lui x18 953391      ====        lui s2, 953391
                                                  30'd    1033    : data = 32'h    B0720593    ;    //    addi x11 x4 -1273      ====        addi a1, tp, -1273
                                                  30'd    1034    : data = 32'h    50E82393    ;    //    slti x7 x16 1294      ====        slti t2, a6, 1294
                                                  30'd    1035    : data = 32'h    010DEC33    ;    //    or x24 x27 x16      ====        or s8, s11, a6
                                                  30'd    1036    : data = 32'h    01BB1B33    ;    //    sll x22 x22 x27      ====        sll s6, s6, s11
                                                  30'd    1037    : data = 32'h    401F0FB3    ;    //    sub x31 x30 x1      ====        sub t6, t5, ra
                                                  30'd    1038    : data = 32'h    F000A713    ;    //    slti x14 x1 -256      ====        slti a4, ra, -256
                                                  30'd    1039    : data = 32'h    01DC1013    ;    //    slli x0 x24 29      ====        slli zero, s8, 29
                                                  30'd    1040    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1041    : data = 32'h    41B155B3    ;    //    sra x11 x2 x27      ====        sra a1, sp, s11
                                                  30'd    1042    : data = 32'h    018B1AB3    ;    //    sll x21 x22 x24      ====        sll s5, s6, s8
                                                  30'd    1043    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1044    : data = 32'h    167CC8B7    ;    //    lui x17 92108      ====        lui a7, 92108
                                                  30'd    1045    : data = 32'h    24D7DC37    ;    //    lui x24 150909      ====        lui s8, 150909
                                                  30'd    1046    : data = 32'h    4018D1B3    ;    //    sra x3 x17 x1      ====        sra gp, a7, ra
                                                  30'd    1047    : data = 32'h    3DDCF317    ;    //    auipc x6 253391      ====        auipc t1, 253391
                                                  30'd    1048    : data = 32'h    F8647593    ;    //    andi x11 x8 -122      ====        andi a1, s0, -122
                                                  30'd    1049    : data = 32'h    6F534693    ;    //    xori x13 x6 1781      ====        xori a3, t1, 1781
                                                  30'd    1050    : data = 32'h    018619B3    ;    //    sll x19 x12 x24      ====        sll s3, a2, s8
                                                  30'd    1051    : data = 32'h    005631B3    ;    //    sltu x3 x12 x5      ====        sltu gp, a2, t0
                                                  30'd    1052    : data = 32'h    4173D313    ;    //    srai x6 x7 23      ====        srai t1, t2, 23
                                                  30'd    1053    : data = 32'h    4B3EDCB7    ;    //    lui x25 308205      ====        lui s9, 308205
                                                  30'd    1054    : data = 32'h    01929A33    ;    //    sll x20 x5 x25      ====        sll s4, t0, s9
                                                  30'd    1055    : data = 32'h    009D5593    ;    //    srli x11 x26 9      ====        srli a1, s10, 9
                                                  30'd    1056    : data = 32'h    408BDB33    ;    //    sra x22 x23 x8      ====        sra s6, s7, s0
                                                  30'd    1057    : data = 32'h    CD168993    ;    //    addi x19 x13 -815      ====        addi s3, a3, -815
                                                  30'd    1058    : data = 32'h    72B9EC13    ;    //    ori x24 x19 1835      ====        ori s8, s3, 1835
                                                  30'd    1059    : data = 32'h    8901BB13    ;    //    sltiu x22 x3 -1904      ====        sltiu s6, gp, -1904
                                                  30'd    1060    : data = 32'h    00AF52B3    ;    //    srl x5 x30 x10      ====        srl t0, t5, a0
                                                  30'd    1061    : data = 32'h    01008FB3    ;    //    add x31 x1 x16      ====        add t6, ra, a6
                                                  30'd    1062    : data = 32'h    48222A93    ;    //    slti x21 x4 1154      ====        slti s5, tp, 1154
                                                  30'd    1063    : data = 32'h    01A1D833    ;    //    srl x16 x3 x26      ====        srl a6, gp, s10
                                                  30'd    1064    : data = 32'h    BA925737    ;    //    lui x14 764197      ====        lui a4, 764197
                                                  30'd    1065    : data = 32'h    96E58613    ;    //    addi x12 x11 -1682      ====        addi a2, a1, -1682
                                                  30'd    1066    : data = 32'h    00E36BB3    ;    //    or x23 x6 x14      ====        or s7, t1, a4
                                                  30'd    1067    : data = 32'h    00FBD493    ;    //    srli x9 x23 15      ====        srli s1, s7, 15
                                                  30'd    1068    : data = 32'h    8593C913    ;    //    xori x18 x7 -1959      ====        xori s2, t2, -1959
                                                  30'd    1069    : data = 32'h    00C194B3    ;    //    sll x9 x3 x12      ====        sll s1, gp, a2
                                                  30'd    1070    : data = 32'h    C9774797    ;    //    auipc x15 825204      ====        auipc a5, 825204
                                                  30'd    1071    : data = 32'h    046C7117    ;    //    auipc x2 18119      ====        auipc sp, 18119
                                                  30'd    1072    : data = 32'h    001E1013    ;    //    slli x0 x28 1      ====        slli zero, t3, 1
                                                  30'd    1073    : data = 32'h    42782D13    ;    //    slti x26 x16 1063      ====        slti s10, a6, 1063
                                                  30'd    1074    : data = 32'h    006028B3    ;    //    slt x17 x0 x6      ====        slt a7, zero, t1
                                                  30'd    1075    : data = 32'h    05E70013    ;    //    addi x0 x14 94      ====        addi zero, a4, 94
                                                  30'd    1076    : data = 32'h    8C872D13    ;    //    slti x26 x14 -1848      ====        slti s10, a4, -1848
                                                  30'd    1077    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1078    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1079    : data = 32'h    CED52437    ;    //    lui x8 847186      ====        lui s0, 847186
                                                  30'd    1080    : data = 32'h    00DA2AB3    ;    //    slt x21 x20 x13      ====        slt s5, s4, a3
                                                  30'd    1081    : data = 32'h    00A57A33    ;    //    and x20 x10 x10      ====        and s4, a0, a0
                                                  30'd    1082    : data = 32'h    01B35E33    ;    //    srl x28 x6 x27      ====        srl t3, t1, s11
                                                  30'd    1083    : data = 32'h    01B239B3    ;    //    sltu x19 x4 x27      ====        sltu s3, tp, s11
                                                  30'd    1084    : data = 32'h    0061D2B3    ;    //    srl x5 x3 x6      ====        srl t0, gp, t1
                                                  30'd    1085    : data = 32'h    90510313    ;    //    addi x6 x2 -1787      ====        addi t1, sp, -1787
                                                  30'd    1086    : data = 32'h    0107DB13    ;    //    srli x22 x15 16      ====        srli s6, a5, 16
                                                  30'd    1087    : data = 32'h    019DF7B3    ;    //    and x15 x27 x25      ====        and a5, s11, s9
                                                  30'd    1088    : data = 32'h    005017B3    ;    //    sll x15 x0 x5      ====        sll a5, zero, t0
                                                  30'd    1089    : data = 32'h    012B9333    ;    //    sll x6 x23 x18      ====        sll t1, s7, s2
                                                  30'd    1090    : data = 32'h    008C44B3    ;    //    xor x9 x24 x8      ====        xor s1, s8, s0
                                                  30'd    1091    : data = 32'h    01741293    ;    //    slli x5 x8 23      ====        slli t0, s0, 23
                                                  30'd    1092    : data = 32'h    00970133    ;    //    add x2 x14 x9      ====        add sp, a4, s1
                                                  30'd    1093    : data = 32'h    418208B3    ;    //    sub x17 x4 x24      ====        sub a7, tp, s8
                                                  30'd    1094    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1095    : data = 32'h    416FD2B3    ;    //    sra x5 x31 x22      ====        sra t0, t6, s6
                                                  30'd    1096    : data = 32'h    33360293    ;    //    addi x5 x12 819      ====        addi t0, a2, 819
                                                  30'd    1097    : data = 32'h    C2EB4697    ;    //    auipc x13 798388      ====        auipc a3, 798388
                                                  30'd    1098    : data = 32'h    016FD033    ;    //    srl x0 x31 x22      ====        srl zero, t6, s6
                                                  30'd    1099    : data = 32'h    008FDCB3    ;    //    srl x25 x31 x8      ====        srl s9, t6, s0
                                                  30'd    1100    : data = 32'h    00258EB3    ;    //    add x29 x11 x2      ====        add t4, a1, sp
                                                  30'd    1101    : data = 32'h    01C98933    ;    //    add x18 x19 x28      ====        add s2, s3, t3
                                                  30'd    1102    : data = 32'h    00985C13    ;    //    srli x24 x16 9      ====        srli s8, a6, 9
                                                  30'd    1103    : data = 32'h    0A35A293    ;    //    slti x5 x11 163      ====        slti t0, a1, 163
                                                  30'd    1104    : data = 32'h    01DADE33    ;    //    srl x28 x21 x29      ====        srl t3, s5, t4
                                                  30'd    1105    : data = 32'h    914EEE93    ;    //    ori x29 x29 -1772      ====        ori t4, t4, -1772
                                                  30'd    1106    : data = 32'h    3D540B93    ;    //    addi x23 x8 981      ====        addi s7, s0, 981
                                                  30'd    1107    : data = 32'h    5F56FB13    ;    //    andi x22 x13 1525      ====        andi s6, a3, 1525
                                                  30'd    1108    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1109    : data = 32'h    00195A13    ;    //    srli x20 x18 1      ====        srli s4, s2, 1
                                                  30'd    1110    : data = 32'h    FF0FEE93    ;    //    ori x29 x31 -16      ====        ori t4, t6, -16
                                                  30'd    1111    : data = 32'h    13B4F393    ;    //    andi x7 x9 315      ====        andi t2, s1, 315
                                                  30'd    1112    : data = 32'h    000EC933    ;    //    xor x18 x29 x0      ====        xor s2, t4, zero
                                                  30'd    1113    : data = 32'h    BBCF3097    ;    //    auipc x1 769267      ====        auipc ra, 769267
                                                  30'd    1114    : data = 32'h    41C159B3    ;    //    sra x19 x2 x28      ====        sra s3, sp, t3
                                                  30'd    1115    : data = 32'h    0026DB93    ;    //    srli x23 x13 2      ====        srli s7, a3, 2
                                                  30'd    1116    : data = 32'h    C314C313    ;    //    xori x6 x9 -975      ====        xori t1, s1, -975
                                                  30'd    1117    : data = 32'h    8EC04193    ;    //    xori x3 x0 -1812      ====        xori gp, zero, -1812
                                                  30'd    1118    : data = 32'h    41D6D193    ;    //    srai x3 x13 29      ====        srai gp, a3, 29
                                                  30'd    1119    : data = 32'h    00A71FB3    ;    //    sll x31 x14 x10      ====        sll t6, a4, a0
                                                  30'd    1120    : data = 32'h    01A53CB3    ;    //    sltu x25 x10 x26      ====        sltu s9, a0, s10
                                                  30'd    1121    : data = 32'h    360BEE13    ;    //    ori x28 x23 864      ====        ori t3, s7, 864
                                                  30'd    1122    : data = 32'h    41CDD933    ;    //    sra x18 x27 x28      ====        sra s2, s11, t3
                                                  30'd    1123    : data = 32'h    DC42AA13    ;    //    slti x20 x5 -572      ====        slti s4, t0, -572
                                                  30'd    1124    : data = 32'h    33F1FA37    ;    //    lui x20 212767      ====        lui s4, 212767
                                                  30'd    1125    : data = 32'h    D55ECB93    ;    //    xori x23 x29 -683      ====        xori s7, t4, -683
                                                  30'd    1126    : data = 32'h    AC2AB893    ;    //    sltiu x17 x21 -1342      ====        sltiu a7, s5, -1342
                                                  30'd    1127    : data = 32'h    A5D23313    ;    //    sltiu x6 x4 -1443      ====        sltiu t1, tp, -1443
                                                  30'd    1128    : data = 32'h    010F0A33    ;    //    add x20 x30 x16      ====        add s4, t5, a6
                                                  30'd    1129    : data = 32'h    007148B3    ;    //    xor x17 x2 x7      ====        xor a7, sp, t2
                                                  30'd    1130    : data = 32'h    F50FE993    ;    //    ori x19 x31 -176      ====        ori s3, t6, -176
                                                  30'd    1131    : data = 32'h    F7E6EC13    ;    //    ori x24 x13 -130      ====        ori s8, a3, -130
                                                  30'd    1132    : data = 32'h    404252B3    ;    //    sra x5 x4 x4      ====        sra t0, tp, tp
                                                  30'd    1133    : data = 32'h    C9331497    ;    //    auipc x9 824113      ====        auipc s1, 824113
                                                  30'd    1134    : data = 32'h    88D37A93    ;    //    andi x21 x6 -1907      ====        andi s5, t1, -1907
                                                  30'd    1135    : data = 32'h    01F51D13    ;    //    slli x26 x10 31      ====        slli s10, a0, 31
                                                  30'd    1136    : data = 32'h    01EB1E33    ;    //    sll x28 x22 x30      ====        sll t3, s6, t5
                                                  30'd    1137    : data = 32'h    4CAE8D93    ;    //    addi x27 x29 1226      ====        addi s11, t4, 1226
                                                  30'd    1138    : data = 32'h    405855B3    ;    //    sra x11 x16 x5      ====        sra a1, a6, t0
                                                  30'd    1139    : data = 32'h    00D22133    ;    //    slt x2 x4 x13      ====        slt sp, tp, a3
                                                  30'd    1140    : data = 32'h    013BA633    ;    //    slt x12 x23 x19      ====        slt a2, s7, s3
                                                  30'd    1141    : data = 32'h    B48CDE97    ;    //    auipc x29 739533      ====        auipc t4, 739533
                                                  30'd    1142    : data = 32'h    0086CCB3    ;    //    xor x25 x13 x8      ====        xor s9, a3, s0
                                                  30'd    1143    : data = 32'h    415D02B3    ;    //    sub x5 x26 x21      ====        sub t0, s10, s5
                                                  30'd    1144    : data = 32'h    41D75D13    ;    //    srai x26 x14 29      ====        srai s10, a4, 29
                                                  30'd    1145    : data = 32'h    40A88C33    ;    //    sub x24 x17 x10      ====        sub s8, a7, a0
                                                  30'd    1146    : data = 32'h    01B51913    ;    //    slli x18 x10 27      ====        slli s2, a0, 27
                                                  30'd    1147    : data = 32'h    479A3713    ;    //    sltiu x14 x20 1145      ====        sltiu a4, s4, 1145
                                                  30'd    1148    : data = 32'h    AC5E7093    ;    //    andi x1 x28 -1339      ====        andi ra, t3, -1339
                                                  30'd    1149    : data = 32'h    00B8BFB3    ;    //    sltu x31 x17 x11      ====        sltu t6, a7, a1
                                                  30'd    1150    : data = 32'h    2230B293    ;    //    sltiu x5 x1 547      ====        sltiu t0, ra, 547
                                                  30'd    1151    : data = 32'h    01991193    ;    //    slli x3 x18 25      ====        slli gp, s2, 25
                                                  30'd    1152    : data = 32'h    01AE8DB3    ;    //    add x27 x29 x26      ====        add s11, t4, s10
                                                  30'd    1153    : data = 32'h    3E1E4913    ;    //    xori x18 x28 993      ====        xori s2, t3, 993
                                                  30'd    1154    : data = 32'h    9232F413    ;    //    andi x8 x5 -1757      ====        andi s0, t0, -1757
                                                  30'd    1155    : data = 32'h    4137D9B3    ;    //    sra x19 x15 x19      ====        sra s3, a5, s3
                                                  30'd    1156    : data = 32'h    B645F393    ;    //    andi x7 x11 -1180      ====        andi t2, a1, -1180
                                                  30'd    1157    : data = 32'h    0EAC7C17    ;    //    auipc x24 60103      ====        auipc s8, 60103
                                                  30'd    1158    : data = 32'h    013D89B3    ;    //    add x19 x27 x19      ====        add s3, s11, s3
                                                  30'd    1159    : data = 32'h    00FA71B3    ;    //    and x3 x20 x15      ====        and gp, s4, a5
                                                  30'd    1160    : data = 32'h    296B0793    ;    //    addi x15 x22 662      ====        addi a5, s6, 662
                                                  30'd    1161    : data = 32'h    41285E33    ;    //    sra x28 x16 x18      ====        sra t3, a6, s2
                                                  30'd    1162    : data = 32'h    D5F46D93    ;    //    ori x27 x8 -673      ====        ori s11, s0, -673
                                                  30'd    1163    : data = 32'h    00874AB3    ;    //    xor x21 x14 x8      ====        xor s5, a4, s0
                                                  30'd    1164    : data = 32'h    016A73B3    ;    //    and x7 x20 x22      ====        and t2, s4, s6
                                                  30'd    1165    : data = 32'h    35F8E917    ;    //    auipc x18 221070      ====        auipc s2, 221070
                                                  30'd    1166    : data = 32'h    4052D733    ;    //    sra x14 x5 x5      ====        sra a4, t0, t0
                                                  30'd    1167    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1168    : data = 32'h    011F6FB3    ;    //    or x31 x30 x17      ====        or t6, t5, a7
                                                  30'd    1169    : data = 32'h    0025E9B3    ;    //    or x19 x11 x2      ====        or s3, a1, sp
                                                  30'd    1170    : data = 32'h    007D9113    ;    //    slli x2 x27 7      ====        slli sp, s11, 7
                                                  30'd    1171    : data = 32'h    01515A93    ;    //    srli x21 x2 21      ====        srli s5, sp, 21
                                                  30'd    1172    : data = 32'h    00DD08B3    ;    //    add x17 x26 x13      ====        add a7, s10, a3
                                                  30'd    1173    : data = 32'h    009DFCB3    ;    //    and x25 x27 x9      ====        and s9, s11, s1
                                                  30'd    1174    : data = 32'h    00F6D5B3    ;    //    srl x11 x13 x15      ====        srl a1, a3, a5
                                                  30'd    1175    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1176    : data = 32'h    406F80B3    ;    //    sub x1 x31 x6      ====        sub ra, t6, t1
                                                  30'd    1177    : data = 32'h    C17CBF93    ;    //    sltiu x31 x25 -1001      ====        sltiu t6, s9, -1001
                                                  30'd    1178    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1179    : data = 32'h    01BC1493    ;    //    slli x9 x24 27      ====        slli s1, s8, 27
                                                  30'd    1180    : data = 32'h    00125B93    ;    //    srli x23 x4 1      ====        srli s7, tp, 1
                                                  30'd    1181    : data = 32'h    40555F93    ;    //    srai x31 x10 5      ====        srai t6, a0, 5
                                                  30'd    1182    : data = 32'h    41980EB3    ;    //    sub x29 x16 x25      ====        sub t4, a6, s9
                                                  30'd    1183    : data = 32'h    4ABC8A13    ;    //    addi x20 x25 1195      ====        addi s4, s9, 1195
                                                  30'd    1184    : data = 32'h    181D2C13    ;    //    slti x24 x26 385      ====        slti s8, s10, 385
                                                  30'd    1185    : data = 32'h    008FADB3    ;    //    slt x27 x31 x8      ====        slt s11, t6, s0
                                                  30'd    1186    : data = 32'h    0015A1B3    ;    //    slt x3 x11 x1      ====        slt gp, a1, ra
                                                  30'd    1187    : data = 32'h    00BB4C33    ;    //    xor x24 x22 x11      ====        xor s8, s6, a1
                                                  30'd    1188    : data = 32'h    01A55593    ;    //    srli x11 x10 26      ====        srli a1, a0, 26
                                                  30'd    1189    : data = 32'h    59806D93    ;    //    ori x27 x0 1432      ====        ori s11, zero, 1432
                                                  30'd    1190    : data = 32'h    0011E2B3    ;    //    or x5 x3 x1      ====        or t0, gp, ra
                                                  30'd    1191    : data = 32'h    5EC7D317    ;    //    auipc x6 388221      ====        auipc t1, 388221
                                                  30'd    1192    : data = 32'h    56910E37    ;    //    lui x28 354576      ====        lui t3, 354576
                                                  30'd    1193    : data = 32'h    0108B5B3    ;    //    sltu x11 x17 x16      ====        sltu a1, a7, a6
                                                  30'd    1194    : data = 32'h    017D1193    ;    //    slli x3 x26 23      ====        slli gp, s10, 23
                                                  30'd    1195    : data = 32'h    001B75B3    ;    //    and x11 x22 x1      ====        and a1, s6, ra
                                                  30'd    1196    : data = 32'h    0006D0B3    ;    //    srl x1 x13 x0      ====        srl ra, a3, zero
                                                  30'd    1197    : data = 32'h    367D6293    ;    //    ori x5 x26 871      ====        ori t0, s10, 871
                                                  30'd    1198    : data = 32'h    C486E017    ;    //    auipc x0 804974      ====        auipc zero, 804974
                                                  30'd    1199    : data = 32'h    01C1D1B3    ;    //    srl x3 x3 x28      ====        srl gp, gp, t3
                                                  30'd    1200    : data = 32'h    EB2A0DB7    ;    //    lui x27 963232      ====        lui s11, 963232
                                                  30'd    1201    : data = 32'h    015352B3    ;    //    srl x5 x6 x21      ====        srl t0, t1, s5
                                                  30'd    1202    : data = 32'h    99783793    ;    //    sltiu x15 x16 -1641      ====        sltiu a5, a6, -1641
                                                  30'd    1203    : data = 32'h    407504B3    ;    //    sub x9 x10 x7      ====        sub s1, a0, t2
                                                  30'd    1204    : data = 32'h    01F00D33    ;    //    add x26 x0 x31      ====        add s10, zero, t6
                                                  30'd    1205    : data = 32'h    0166DE13    ;    //    srli x28 x13 22      ====        srli t3, a3, 22
                                                  30'd    1206    : data = 32'h    8F1E3897    ;    //    auipc x17 586211      ====        auipc a7, 586211
                                                  30'd    1207    : data = 32'h    008156B3    ;    //    srl x13 x2 x8      ====        srl a3, sp, s0
                                                  30'd    1208    : data = 32'h    005A5893    ;    //    srli x17 x20 5      ====        srli a7, s4, 5
                                                  30'd    1209    : data = 32'h    40B908B3    ;    //    sub x17 x18 x11      ====        sub a7, s2, a1
                                                  30'd    1210    : data = 32'h    0168B933    ;    //    sltu x18 x17 x22      ====        sltu s2, a7, s6
                                                  30'd    1211    : data = 32'h    01C71013    ;    //    slli x0 x14 28      ====        slli zero, a4, 28
                                                  30'd    1212    : data = 32'h    0183A033    ;    //    slt x0 x7 x24      ====        slt zero, t2, s8
                                                  30'd    1213    : data = 32'h    416E5C93    ;    //    srai x25 x28 22      ====        srai s9, t3, 22
                                                  30'd    1214    : data = 32'h    008D8933    ;    //    add x18 x27 x8      ====        add s2, s11, s0
                                                  30'd    1215    : data = 32'h    1CD50B97    ;    //    auipc x23 118096      ====        auipc s7, 118096
                                                  30'd    1216    : data = 32'h    01781C33    ;    //    sll x24 x16 x23      ====        sll s8, a6, s7
                                                  30'd    1217    : data = 32'h    41015133    ;    //    sra x2 x2 x16      ====        sra sp, sp, a6
                                                  30'd    1218    : data = 32'h    00739F93    ;    //    slli x31 x7 7      ====        slli t6, t2, 7
                                                  30'd    1219    : data = 32'h    00979D13    ;    //    slli x26 x15 9      ====        slli s10, a5, 9
                                                  30'd    1220    : data = 32'h    013AB0B3    ;    //    sltu x1 x21 x19      ====        sltu ra, s5, s3
                                                  30'd    1221    : data = 32'h    000A5CB3    ;    //    srl x25 x20 x0      ====        srl s9, s4, zero
                                                  30'd    1222    : data = 32'h    4E6F4A17    ;    //    auipc x20 321268      ====        auipc s4, 321268
                                                  30'd    1223    : data = 32'h    00978733    ;    //    add x14 x15 x9      ====        add a4, a5, s1
                                                  30'd    1224    : data = 32'h    D9FFDA37    ;    //    lui x20 892925      ====        lui s4, 892925
                                                  30'd    1225    : data = 32'h    41F3DAB3    ;    //    sra x21 x7 x31      ====        sra s5, t2, t6
                                                  30'd    1226    : data = 32'h    01DEA333    ;    //    slt x6 x29 x29      ====        slt t1, t4, t4
                                                  30'd    1227    : data = 32'h    01245E93    ;    //    srli x29 x8 18      ====        srli t4, s0, 18
                                                  30'd    1228    : data = 32'h    01F03733    ;    //    sltu x14 x0 x31      ====        sltu a4, zero, t6
                                                  30'd    1229    : data = 32'h    01E4EDB3    ;    //    or x27 x9 x30      ====        or s11, s1, t5
                                                  30'd    1230    : data = 32'h    010AD593    ;    //    srli x11 x21 16      ====        srli a1, s5, 16
                                                  30'd    1231    : data = 32'h    006D1613    ;    //    slli x12 x26 6      ====        slli a2, s10, 6
                                                  30'd    1232    : data = 32'h    E067B013    ;    //    sltiu x0 x15 -506      ====        sltiu zero, a5, -506
                                                  30'd    1233    : data = 32'h    0094A6B3    ;    //    slt x13 x9 x9      ====        slt a3, s1, s1
                                                  30'd    1234    : data = 32'h    3DA83593    ;    //    sltiu x11 x16 986      ====        sltiu a1, a6, 986
                                                  30'd    1235    : data = 32'h    00803933    ;    //    sltu x18 x0 x8      ====        sltu s2, zero, s0
                                                  30'd    1236    : data = 32'h    00E8BBB3    ;    //    sltu x23 x17 x14      ====        sltu s7, a7, a4
                                                  30'd    1237    : data = 32'h    D9607E93    ;    //    andi x29 x0 -618      ====        andi t4, zero, -618
                                                  30'd    1238    : data = 32'h    4A1B6817    ;    //    auipc x16 303542      ====        auipc a6, 303542
                                                  30'd    1239    : data = 32'h    3CD77593    ;    //    andi x11 x14 973      ====        andi a1, a4, 973
                                                  30'd    1240    : data = 32'h    2B168093    ;    //    addi x1 x13 689      ====        addi ra, a3, 689
                                                  30'd    1241    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1242    : data = 32'h    0076F3B3    ;    //    and x7 x13 x7      ====        and t2, a3, t2
                                                  30'd    1243    : data = 32'h    ED930A13    ;    //    addi x20 x6 -295      ====        addi s4, t1, -295
                                                  30'd    1244    : data = 32'h    68E0FB13    ;    //    andi x22 x1 1678      ====        andi s6, ra, 1678
                                                  30'd    1245    : data = 32'h    F88E7293    ;    //    andi x5 x28 -120      ====        andi t0, t3, -120
                                                  30'd    1246    : data = 32'h    D4DF3413    ;    //    sltiu x8 x30 -691      ====        sltiu s0, t5, -691
                                                  30'd    1247    : data = 32'h    AC76D8B7    ;    //    lui x17 706413      ====        lui a7, 706413
                                                  30'd    1248    : data = 32'h    0182A333    ;    //    slt x6 x5 x24      ====        slt t1, t0, s8
                                                  30'd    1249    : data = 32'h    094F2713    ;    //    slti x14 x30 148      ====        slti a4, t5, 148
                                                  30'd    1250    : data = 32'h    01F30333    ;    //    add x6 x6 x31      ====        add t1, t1, t6
                                                  30'd    1251    : data = 32'h    34F00093    ;    //    addi x1 x0 847      ====        addi ra, zero, 847
                                                  30'd    1252    : data = 32'h    0144EA33    ;    //    or x20 x9 x20      ====        or s4, s1, s4
                                                  30'd    1253    : data = 32'h    01423033    ;    //    sltu x0 x4 x20      ====        sltu zero, tp, s4
                                                  30'd    1254    : data = 32'h    5799F313    ;    //    andi x6 x19 1401      ====        andi t1, s3, 1401
                                                  30'd    1255    : data = 32'h    D003B593    ;    //    sltiu x11 x7 -768      ====        sltiu a1, t2, -768
                                                  30'd    1256    : data = 32'h    3018FB93    ;    //    andi x23 x17 769      ====        andi s7, a7, 769
                                                  30'd    1257    : data = 32'h    019BC833    ;    //    xor x16 x23 x25      ====        xor a6, s7, s9
                                                  30'd    1258    : data = 32'h    009FC433    ;    //    xor x8 x31 x9      ====        xor s0, t6, s1
                                                  30'd    1259    : data = 32'h    01EEE3B3    ;    //    or x7 x29 x30      ====        or t2, t4, t5
                                                  30'd    1260    : data = 32'h    00A6BE33    ;    //    sltu x28 x13 x10      ====        sltu t3, a3, a0
                                                  30'd    1261    : data = 32'h    01DB2133    ;    //    slt x2 x22 x29      ====        slt sp, s6, t4
                                                  30'd    1262    : data = 32'h    00F5B033    ;    //    sltu x0 x11 x15      ====        sltu zero, a1, a5
                                                  30'd    1263    : data = 32'h    00071A33    ;    //    sll x20 x14 x0      ====        sll s4, a4, zero
                                                  30'd    1264    : data = 32'h    000F9D13    ;    //    slli x26 x31 0      ====        slli s10, t6, 0
                                                  30'd    1265    : data = 32'h    00E9AAB3    ;    //    slt x21 x19 x14      ====        slt s5, s3, a4
                                                  30'd    1266    : data = 32'h    97B37C13    ;    //    andi x24 x6 -1669      ====        andi s8, t1, -1669
                                                  30'd    1267    : data = 32'h    90FBF413    ;    //    andi x8 x23 -1777      ====        andi s0, s7, -1777
                                                  30'd    1268    : data = 32'h    415B5293    ;    //    srai x5 x22 21      ====        srai t0, s6, 21
                                                  30'd    1269    : data = 32'h    A5C032B7    ;    //    lui x5 678915      ====        lui t0, 678915
                                                  30'd    1270    : data = 32'h    41BF8633    ;    //    sub x12 x31 x27      ====        sub a2, t6, s11
                                                  30'd    1271    : data = 32'h    3EB76893    ;    //    ori x17 x14 1003      ====        ori a7, a4, 1003
                                                  30'd    1272    : data = 32'h    01303C33    ;    //    sltu x24 x0 x19      ====        sltu s8, zero, s3
                                                  30'd    1273    : data = 32'h    40D8C593    ;    //    xori x11 x17 1037      ====        xori a1, a7, 1037
                                                  30'd    1274    : data = 32'h    00D4EDB3    ;    //    or x27 x9 x13      ====        or s11, s1, a3
                                                  30'd    1275    : data = 32'h    D3D78993    ;    //    addi x19 x15 -707      ====        addi s3, a5, -707
                                                  30'd    1276    : data = 32'h    0171D993    ;    //    srli x19 x3 23      ====        srli s3, gp, 23
                                                  30'd    1277    : data = 32'h    014C27B3    ;    //    slt x15 x24 x20      ====        slt a5, s8, s4
                                                  30'd    1278    : data = 32'h    305D0613    ;    //    addi x12 x26 773      ====        addi a2, s10, 773
                                                  30'd    1279    : data = 32'h    39B17793    ;    //    andi x15 x2 923      ====        andi a5, sp, 923
                                                  30'd    1280    : data = 32'h    2A032197    ;    //    auipc x3 172082      ====        auipc gp, 172082
                                                  30'd    1281    : data = 32'h    01D9B733    ;    //    sltu x14 x19 x29      ====        sltu a4, s3, t4
                                                  30'd    1282    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1283    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1284    : data = 32'h    52C76593    ;    //    ori x11 x14 1324      ====        ori a1, a4, 1324
                                                  30'd    1285    : data = 32'h    2D3D2E13    ;    //    slti x28 x26 723      ====        slti t3, s10, 723
                                                  30'd    1286    : data = 32'h    40C0D033    ;    //    sra x0 x1 x12      ====        sra zero, ra, a2
                                                  30'd    1287    : data = 32'h    00E637B3    ;    //    sltu x15 x12 x14      ====        sltu a5, a2, a4
                                                  30'd    1288    : data = 32'h    0116F9B3    ;    //    and x19 x13 x17      ====        and s3, a3, a7
                                                  30'd    1289    : data = 32'h    0115DD33    ;    //    srl x26 x11 x17      ====        srl s10, a1, a7
                                                  30'd    1290    : data = 32'h    EC2ABB13    ;    //    sltiu x22 x21 -318      ====        sltiu s6, s5, -318
                                                  30'd    1291    : data = 32'h    24B93793    ;    //    sltiu x15 x18 587      ====        sltiu a5, s2, 587
                                                  30'd    1292    : data = 32'h    41898413    ;    //    addi x8 x19 1048      ====        addi s0, s3, 1048
                                                  30'd    1293    : data = 32'h    01A2BE33    ;    //    sltu x28 x5 x26      ====        sltu t3, t0, s10
                                                  30'd    1294    : data = 32'h    41DB5493    ;    //    srai x9 x22 29      ====        srai s1, s6, 29
                                                  30'd    1295    : data = 32'h    01C5ABB3    ;    //    slt x23 x11 x28      ====        slt s7, a1, t3
                                                  30'd    1296    : data = 32'h    00D033B3    ;    //    sltu x7 x0 x13      ====        sltu t2, zero, a3
                                                  30'd    1297    : data = 32'h    0192DF93    ;    //    srli x31 x5 25      ====        srli t6, t0, 25
                                                  30'd    1298    : data = 32'h    98CA7813    ;    //    andi x16 x20 -1652      ====        andi a6, s4, -1652
                                                  30'd    1299    : data = 32'h    01185B33    ;    //    srl x22 x16 x17      ====        srl s6, a6, a7
                                                  30'd    1300    : data = 32'h    008E64B3    ;    //    or x9 x28 x8      ====        or s1, t3, s0
                                                  30'd    1301    : data = 32'h    D0134713    ;    //    xori x14 x6 -767      ====        xori a4, t1, -767
                                                  30'd    1302    : data = 32'h    018C2333    ;    //    slt x6 x24 x24      ====        slt t1, s8, s8
                                                  30'd    1303    : data = 32'h    5C5D4893    ;    //    xori x17 x26 1477      ====        xori a7, s10, 1477
                                                  30'd    1304    : data = 32'h    C8AAC793    ;    //    xori x15 x21 -886      ====        xori a5, s5, -886
                                                  30'd    1305    : data = 32'h    D92A0693    ;    //    addi x13 x20 -622      ====        addi a3, s4, -622
                                                  30'd    1306    : data = 32'h    000E4933    ;    //    xor x18 x28 x0      ====        xor s2, t3, zero
                                                  30'd    1307    : data = 32'h    C5D48313    ;    //    addi x6 x9 -931      ====        addi t1, s1, -931
                                                  30'd    1308    : data = 32'h    4034DFB3    ;    //    sra x31 x9 x3      ====        sra t6, s1, gp
                                                  30'd    1309    : data = 32'h    0005C433    ;    //    xor x8 x11 x0      ====        xor s0, a1, zero
                                                  30'd    1310    : data = 32'h    7E513B13    ;    //    sltiu x22 x2 2021      ====        sltiu s6, sp, 2021
                                                  30'd    1311    : data = 32'h    01B79733    ;    //    sll x14 x15 x27      ====        sll a4, a5, s11
                                                  30'd    1312    : data = 32'h    4163D713    ;    //    srai x14 x7 22      ====        srai a4, t2, 22
                                                  30'd    1313    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1314    : data = 32'h    B7FD4E37    ;    //    lui x28 753620      ====        lui t3, 753620
                                                  30'd    1315    : data = 32'h    41718633    ;    //    sub x12 x3 x23      ====        sub a2, gp, s7
                                                  30'd    1316    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1317    : data = 32'h    01F94E33    ;    //    xor x28 x18 x31      ====        xor t3, s2, t6
                                                  30'd    1318    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1319    : data = 32'h    00FF4633    ;    //    xor x12 x30 x15      ====        xor a2, t5, a5
                                                  30'd    1320    : data = 32'h    40625B93    ;    //    srai x23 x4 6      ====        srai s7, tp, 6
                                                  30'd    1321    : data = 32'h    41495093    ;    //    srai x1 x18 20      ====        srai ra, s2, 20
                                                  30'd    1322    : data = 32'h    40D05A33    ;    //    sra x20 x0 x13      ====        sra s4, zero, a3
                                                  30'd    1323    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1324    : data = 32'h    EDC5A993    ;    //    slti x19 x11 -292      ====        slti s3, a1, -292
                                                  30'd    1325    : data = 32'h    01D8D113    ;    //    srli x2 x17 29      ====        srli sp, a7, 29
                                                  30'd    1326    : data = 32'h    0163B3B3    ;    //    sltu x7 x7 x22      ====        sltu t2, t2, s6
                                                  30'd    1327    : data = 32'h    8AA92C93    ;    //    slti x25 x18 -1878      ====        slti s9, s2, -1878
                                                  30'd    1328    : data = 32'h    247CC593    ;    //    xori x11 x25 583      ====        xori a1, s9, 583
                                                  30'd    1329    : data = 32'h    0059A1B3    ;    //    slt x3 x19 x5      ====        slt gp, s3, t0
                                                  30'd    1330    : data = 32'h    01635193    ;    //    srli x3 x6 22      ====        srli gp, t1, 22
                                                  30'd    1331    : data = 32'h    55557993    ;    //    andi x19 x10 1365      ====        andi s3, a0, 1365
                                                  30'd    1332    : data = 32'h    A5D94313    ;    //    xori x6 x18 -1443      ====        xori t1, s2, -1443
                                                  30'd    1333    : data = 32'h    41D0DC33    ;    //    sra x24 x1 x29      ====        sra s8, ra, t4
                                                  30'd    1334    : data = 32'h    01A1B7B3    ;    //    sltu x15 x3 x26      ====        sltu a5, gp, s10
                                                  30'd    1335    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1336    : data = 32'h    6FD0BA93    ;    //    sltiu x21 x1 1789      ====        sltiu s5, ra, 1789
                                                  30'd    1337    : data = 32'h    01469E33    ;    //    sll x28 x13 x20      ====        sll t3, a3, s4
                                                  30'd    1338    : data = 32'h    00000693    ;    //    addi x13 x0 0      ====        li a3, 0x0 #start riscv_int_numeric_corner_stream_8
                                                  30'd    1339    : data = 32'h    80000837    ;    //    lui x16 524288      ====        li a6, 0x80000000
                                                  30'd    1340    : data = 32'h    00080813    ;    //    addi x16 x16 0      ====        li a6, 0x80000000
                                                  30'd    1341    : data = 32'h    800009B7    ;    //    lui x19 524288      ====        li s3, 0x80000000
                                                  30'd    1342    : data = 32'h    00098993    ;    //    addi x19 x19 0      ====        li s3, 0x80000000
                                                  30'd    1343    : data = 32'h    6A590EB7    ;    //    lui x29 435600      ====        li t4, 0x6a59005a
                                                  30'd    1344    : data = 32'h    05AE8E93    ;    //    addi x29 x29 90      ====        li t4, 0x6a59005a
                                                  30'd    1345    : data = 32'h    00000193    ;    //    addi x3 x0 0      ====        li gp, 0x0
                                                  30'd    1346    : data = 32'h    00000A13    ;    //    addi x20 x0 0      ====        li s4, 0x0
                                                  30'd    1347    : data = 32'h    FFF00893    ;    //    addi x17 x0 -1      ====        li a7, 0xffffffff
                                                  30'd    1348    : data = 32'h    00000593    ;    //    addi x11 x0 0      ====        li a1, 0x0
                                                  30'd    1349    : data = 32'h    80000D37    ;    //    lui x26 524288      ====        li s10, 0x80000000
                                                  30'd    1350    : data = 32'h    000D0D13    ;    //    addi x26 x26 0      ====        li s10, 0x80000000
                                                  30'd    1351    : data = 32'h    FFF00793    ;    //    addi x15 x0 -1      ====        li a5, 0xffffffff
                                                  30'd    1352    : data = 32'h    2C8A8E97    ;    //    auipc x29 182440      ====        auipc t4, 182440
                                                  30'd    1353    : data = 32'h    41D88EB3    ;    //    sub x29 x17 x29      ====        sub t4, a7, t4
                                                  30'd    1354    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1355    : data = 32'h    B3A58693    ;    //    addi x13 x11 -1222      ====        addi a3, a1, -1222
                                                  30'd    1356    : data = 32'h    413686B3    ;    //    sub x13 x13 x19      ====        sub a3, a3, s3
                                                  30'd    1357    : data = 32'h    00FE87B3    ;    //    add x15 x29 x15      ====        add a5, t4, a5
                                                  30'd    1358    : data = 32'h    6F613837    ;    //    lui x16 456211      ====        lui a6, 456211
                                                  30'd    1359    : data = 32'h    01058A33    ;    //    add x20 x11 x16      ====        add s4, a1, a6
                                                  30'd    1360    : data = 32'h    0394C7B7    ;    //    lui x15 14668      ====        lui a5, 14668
                                                  30'd    1361    : data = 32'h    EEDE9D17    ;    //    auipc x26 978409      ====        auipc s10, 978409
                                                  30'd    1362    : data = 32'h    403587B3    ;    //    sub x15 x11 x3      ====        sub a5, a1, gp
                                                  30'd    1363    : data = 32'h    94980793    ;    //    addi x15 x16 -1719      ====        addi a5, a6, -1719
                                                  30'd    1364    : data = 32'h    40F807B3    ;    //    sub x15 x16 x15      ====        sub a5, a6, a5
                                                  30'd    1365    : data = 32'h    9D43FD17    ;    //    auipc x26 644159      ====        auipc s10, 644159
                                                  30'd    1366    : data = 32'h    286D0D13    ;    //    addi x26 x26 646      ====        addi s10, s10, 646
                                                  30'd    1367    : data = 32'h    1DE80793    ;    //    addi x15 x16 478      ====        addi a5, a6, 478
                                                  30'd    1368    : data = 32'h    96F88193    ;    //    addi x3 x17 -1681      ====        addi gp, a7, -1681
                                                  30'd    1369    : data = 32'h    00398833    ;    //    add x16 x19 x3      ====        add a6, s3, gp
                                                  30'd    1370    : data = 32'h    1800A0EF    ;    //    jal x1 41344      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_8
                                                  30'd    1371    : data = 32'h    353DA093    ;    //    slti x1 x27 851      ====        slti ra, s11, 851
                                                  30'd    1372    : data = 32'h    178BC413    ;    //    xori x8 x23 376      ====        xori s0, s7, 376
                                                  30'd    1373    : data = 32'h    010F6733    ;    //    or x14 x30 x16      ====        or a4, t5, a6
                                                  30'd    1374    : data = 32'h    41873AB7    ;    //    lui x21 268403      ====        lui s5, 268403
                                                  30'd    1375    : data = 32'h    0180B3B3    ;    //    sltu x7 x1 x24      ====        sltu t2, ra, s8
                                                  30'd    1376    : data = 32'h    500A7493    ;    //    andi x9 x20 1280      ====        andi s1, s4, 1280
                                                  30'd    1377    : data = 32'h    0120C733    ;    //    xor x14 x1 x18      ====        xor a4, ra, s2
                                                  30'd    1378    : data = 32'h    41325933    ;    //    sra x18 x4 x19      ====        sra s2, tp, s3
                                                  30'd    1379    : data = 32'h    B9C0E913    ;    //    ori x18 x1 -1124      ====        ori s2, ra, -1124
                                                  30'd    1380    : data = 32'h    011F6DB3    ;    //    or x27 x30 x17      ====        or s11, t5, a7
                                                  30'd    1381    : data = 32'h    40530B33    ;    //    sub x22 x6 x5      ====        sub s6, t1, t0
                                                  30'd    1382    : data = 32'h    97A1E493    ;    //    ori x9 x3 -1670      ====        ori s1, gp, -1670
                                                  30'd    1383    : data = 32'h    01C3B5B3    ;    //    sltu x11 x7 x28      ====        sltu a1, t2, t3
                                                  30'd    1384    : data = 32'h    1C1A2893    ;    //    slti x17 x20 449      ====        slti a7, s4, 449
                                                  30'd    1385    : data = 32'h    238A9437    ;    //    lui x8 145577      ====        lui s0, 145577
                                                  30'd    1386    : data = 32'h    7054A313    ;    //    slti x6 x9 1797      ====        slti t1, s1, 1797
                                                  30'd    1387    : data = 32'h    EDC92E93    ;    //    slti x29 x18 -292      ====        slti t4, s2, -292
                                                  30'd    1388    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1389    : data = 32'h    406BDA33    ;    //    sra x20 x23 x6      ====        sra s4, s7, t1
                                                  30'd    1390    : data = 32'h    0145DE13    ;    //    srli x28 x11 20      ====        srli t3, a1, 20
                                                  30'd    1391    : data = 32'h    47356A13    ;    //    ori x20 x10 1139      ====        ori s4, a0, 1139
                                                  30'd    1392    : data = 32'h    2D11E613    ;    //    ori x12 x3 721      ====        ori a2, gp, 721
                                                  30'd    1393    : data = 32'h    00015433    ;    //    srl x8 x2 x0      ====        srl s0, sp, zero
                                                  30'd    1394    : data = 32'h    009BB5B3    ;    //    sltu x11 x23 x9      ====        sltu a1, s7, s1
                                                  30'd    1395    : data = 32'h    0173CBB3    ;    //    xor x23 x7 x23      ====        xor s7, t2, s7
                                                  30'd    1396    : data = 32'h    41580433    ;    //    sub x8 x16 x21      ====        sub s0, a6, s5
                                                  30'd    1397    : data = 32'h    00D650B3    ;    //    srl x1 x12 x13      ====        srl ra, a2, a3
                                                  30'd    1398    : data = 32'h    011095B3    ;    //    sll x11 x1 x17      ====        sll a1, ra, a7
                                                  30'd    1399    : data = 32'h    00257133    ;    //    and x2 x10 x2      ====        and sp, a0, sp
                                                  30'd    1400    : data = 32'h    3D9A8313    ;    //    addi x6 x21 985      ====        addi t1, s5, 985
                                                  30'd    1401    : data = 32'h    1010B893    ;    //    sltiu x17 x1 257      ====        sltiu a7, ra, 257
                                                  30'd    1402    : data = 32'h    F18213B7    ;    //    lui x7 989217      ====        lui t2, 989217
                                                  30'd    1403    : data = 32'h    91304D93    ;    //    xori x27 x0 -1773      ====        xori s11, zero, -1773
                                                  30'd    1404    : data = 32'h    01D8DA13    ;    //    srli x20 x17 29      ====        srli s4, a7, 29
                                                  30'd    1405    : data = 32'h    40D30833    ;    //    sub x16 x6 x13      ====        sub a6, t1, a3
                                                  30'd    1406    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1407    : data = 32'h    D4BF6293    ;    //    ori x5 x30 -693      ====        ori t0, t5, -693
                                                  30'd    1408    : data = 32'h    40125093    ;    //    srai x1 x4 1      ====        srai ra, tp, 1
                                                  30'd    1409    : data = 32'h    018FD713    ;    //    srli x14 x31 24      ====        srli a4, t6, 24
                                                  30'd    1410    : data = 32'h    013C7433    ;    //    and x8 x24 x19      ====        and s0, s8, s3
                                                  30'd    1411    : data = 32'h    6CD73593    ;    //    sltiu x11 x14 1741      ====        sltiu a1, a4, 1741
                                                  30'd    1412    : data = 32'h    0CA40E97    ;    //    auipc x29 51776      ====        auipc t4, 51776
                                                  30'd    1413    : data = 32'h    00A859B3    ;    //    srl x19 x16 x10      ====        srl s3, a6, a0
                                                  30'd    1414    : data = 32'h    F87A7413    ;    //    andi x8 x20 -121      ====        andi s0, s4, -121
                                                  30'd    1415    : data = 32'h    00CF1093    ;    //    slli x1 x30 12      ====        slli ra, t5, 12
                                                  30'd    1416    : data = 32'h    00E3EDB3    ;    //    or x27 x7 x14      ====        or s11, t2, a4
                                                  30'd    1417    : data = 32'h    01F13C33    ;    //    sltu x24 x2 x31      ====        sltu s8, sp, t6
                                                  30'd    1418    : data = 32'h    41745933    ;    //    sra x18 x8 x23      ====        sra s2, s0, s7
                                                  30'd    1419    : data = 32'h    0173A5B3    ;    //    slt x11 x7 x23      ====        slt a1, t2, s7
                                                  30'd    1420    : data = 32'h    008E6E33    ;    //    or x28 x28 x8      ====        or t3, t3, s0
                                                  30'd    1421    : data = 32'h    706C3013    ;    //    sltiu x0 x24 1798      ====        sltiu zero, s8, 1798
                                                  30'd    1422    : data = 32'h    8262E317    ;    //    auipc x6 534062      ====        auipc t1, 534062
                                                  30'd    1423    : data = 32'h    41EE89B3    ;    //    sub x19 x29 x30      ====        sub s3, t4, t5
                                                  30'd    1424    : data = 32'h    004A9493    ;    //    slli x9 x21 4      ====        slli s1, s5, 4
                                                  30'd    1425    : data = 32'h    005E3BB3    ;    //    sltu x23 x28 x5      ====        sltu s7, t3, t0
                                                  30'd    1426    : data = 32'h    E3EFA897    ;    //    auipc x17 933626      ====        auipc a7, 933626
                                                  30'd    1427    : data = 32'h    1D759AB7    ;    //    lui x21 120665      ====        lui s5, 120665
                                                  30'd    1428    : data = 32'h    09994193    ;    //    xori x3 x18 153      ====        xori gp, s2, 153
                                                  30'd    1429    : data = 32'h    01A21713    ;    //    slli x14 x4 26      ====        slli a4, tp, 26
                                                  30'd    1430    : data = 32'h    000B5913    ;    //    srli x18 x22 0      ====        srli s2, s6, 0
                                                  30'd    1431    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1432    : data = 32'h    C21A4B93    ;    //    xori x23 x20 -991      ====        xori s7, s4, -991
                                                  30'd    1433    : data = 32'h    1309C393    ;    //    xori x7 x19 304      ====        xori t2, s3, 304
                                                  30'd    1434    : data = 32'h    41430833    ;    //    sub x16 x6 x20      ====        sub a6, t1, s4
                                                  30'd    1435    : data = 32'h    410C85B3    ;    //    sub x11 x25 x16      ====        sub a1, s9, a6
                                                  30'd    1436    : data = 32'h    0049A5B3    ;    //    slt x11 x19 x4      ====        slt a1, s3, tp
                                                  30'd    1437    : data = 32'h    9EA54F93    ;    //    xori x31 x10 -1558      ====        xori t6, a0, -1558
                                                  30'd    1438    : data = 32'h    D07CAE13    ;    //    slti x28 x25 -761      ====        slti t3, s9, -761
                                                  30'd    1439    : data = 32'h    6F8E49B7    ;    //    lui x19 456932      ====        lui s3, 456932
                                                  30'd    1440    : data = 32'h    00B7E9B3    ;    //    or x19 x15 x11      ====        or s3, a5, a1
                                                  30'd    1441    : data = 32'h    008EEB33    ;    //    or x22 x29 x8      ====        or s6, t4, s0
                                                  30'd    1442    : data = 32'h    40D302B3    ;    //    sub x5 x6 x13      ====        sub t0, t1, a3
                                                  30'd    1443    : data = 32'h    01408733    ;    //    add x14 x1 x20      ====        add a4, ra, s4
                                                  30'd    1444    : data = 32'h    400A8FB3    ;    //    sub x31 x21 x0      ====        sub t6, s5, zero
                                                  30'd    1445    : data = 32'h    16438413    ;    //    addi x8 x7 356      ====        addi s0, t2, 356
                                                  30'd    1446    : data = 32'h    10C93C93    ;    //    sltiu x25 x18 268      ====        sltiu s9, s2, 268
                                                  30'd    1447    : data = 32'h    412FD193    ;    //    srai x3 x31 18      ====        srai gp, t6, 18
                                                  30'd    1448    : data = 32'h    01310D33    ;    //    add x26 x2 x19      ====        add s10, sp, s3
                                                  30'd    1449    : data = 32'h    01EC9313    ;    //    slli x6 x25 30      ====        slli t1, s9, 30
                                                  30'd    1450    : data = 32'h    01DE0BB3    ;    //    add x23 x28 x29      ====        add s7, t3, t4
                                                  30'd    1451    : data = 32'h    00F13A33    ;    //    sltu x20 x2 x15      ====        sltu s4, sp, a5
                                                  30'd    1452    : data = 32'h    007C21B3    ;    //    slt x3 x24 x7      ====        slt gp, s8, t2
                                                  30'd    1453    : data = 32'h    01CC88B3    ;    //    add x17 x25 x28      ====        add a7, s9, t3
                                                  30'd    1454    : data = 32'h    90F82593    ;    //    slti x11 x16 -1777      ====        slti a1, a6, -1777
                                                  30'd    1455    : data = 32'h    C0076013    ;    //    ori x0 x14 -1024      ====        ori zero, a4, -1024
                                                  30'd    1456    : data = 32'h    01C29C33    ;    //    sll x24 x5 x28      ====        sll s8, t0, t3
                                                  30'd    1457    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1458    : data = 32'h    00B4DB13    ;    //    srli x22 x9 11      ====        srli s6, s1, 11
                                                  30'd    1459    : data = 32'h    01199DB3    ;    //    sll x27 x19 x17      ====        sll s11, s3, a7
                                                  30'd    1460    : data = 32'h    416459B3    ;    //    sra x19 x8 x22      ====        sra s3, s0, s6
                                                  30'd    1461    : data = 32'h    00328AB3    ;    //    add x21 x5 x3      ====        add s5, t0, gp
                                                  30'd    1462    : data = 32'h    60BDA093    ;    //    slti x1 x27 1547      ====        slti ra, s11, 1547
                                                  30'd    1463    : data = 32'h    4F770A13    ;    //    addi x20 x14 1271      ====        addi s4, a4, 1271
                                                  30'd    1464    : data = 32'h    000C93B3    ;    //    sll x7 x25 x0      ====        sll t2, s9, zero
                                                  30'd    1465    : data = 32'h    002AD093    ;    //    srli x1 x21 2      ====        srli ra, s5, 2
                                                  30'd    1466    : data = 32'h    0047F433    ;    //    and x8 x15 x4      ====        and s0, a5, tp
                                                  30'd    1467    : data = 32'h    008484B3    ;    //    add x9 x9 x8      ====        add s1, s1, s0
                                                  30'd    1468    : data = 32'h    00181E33    ;    //    sll x28 x16 x1      ====        sll t3, a6, ra
                                                  30'd    1469    : data = 32'h    B296F193    ;    //    andi x3 x13 -1239      ====        andi gp, a3, -1239
                                                  30'd    1470    : data = 32'h    40055013    ;    //    srai x0 x10 0      ====        srai zero, a0, 0
                                                  30'd    1471    : data = 32'h    0032D793    ;    //    srli x15 x5 3      ====        srli a5, t0, 3
                                                  30'd    1472    : data = 32'h    01D1AE33    ;    //    slt x28 x3 x29      ====        slt t3, gp, t4
                                                  30'd    1473    : data = 32'h    019D1D13    ;    //    slli x26 x26 25      ====        slli s10, s10, 25
                                                  30'd    1474    : data = 32'h    018F05B3    ;    //    add x11 x30 x24      ====        add a1, t5, s8
                                                  30'd    1475    : data = 32'h    415A5833    ;    //    sra x16 x20 x21      ====        sra a6, s4, s5
                                                  30'd    1476    : data = 32'h    000F9113    ;    //    slli x2 x31 0      ====        slli sp, t6, 0
                                                  30'd    1477    : data = 32'h    A7A70C13    ;    //    addi x24 x14 -1414      ====        addi s8, a4, -1414
                                                  30'd    1478    : data = 32'h    011706B3    ;    //    add x13 x14 x17      ====        add a3, a4, a7
                                                  30'd    1479    : data = 32'h    91B1EA13    ;    //    ori x20 x3 -1765      ====        ori s4, gp, -1765
                                                  30'd    1480    : data = 32'h    A9406093    ;    //    ori x1 x0 -1388      ====        ori ra, zero, -1388
                                                  30'd    1481    : data = 32'h    161D4297    ;    //    auipc x5 90580      ====        auipc t0, 90580
                                                  30'd    1482    : data = 32'h    9E1CB193    ;    //    sltiu x3 x25 -1567      ====        sltiu gp, s9, -1567
                                                  30'd    1483    : data = 32'h    013B6DB3    ;    //    or x27 x22 x19      ====        or s11, s6, s3
                                                  30'd    1484    : data = 32'h    97FAA193    ;    //    slti x3 x21 -1665      ====        slti gp, s5, -1665
                                                  30'd    1485    : data = 32'h    4D68B613    ;    //    sltiu x12 x17 1238      ====        sltiu a2, a7, 1238
                                                  30'd    1486    : data = 32'h    00331713    ;    //    slli x14 x6 3      ====        slli a4, t1, 3
                                                  30'd    1487    : data = 32'h    011A8C33    ;    //    add x24 x21 x17      ====        add s8, s5, a7
                                                  30'd    1488    : data = 32'h    011755B3    ;    //    srl x11 x14 x17      ====        srl a1, a4, a7
                                                  30'd    1489    : data = 32'h    00B65C13    ;    //    srli x24 x12 11      ====        srli s8, a2, 11
                                                  30'd    1490    : data = 32'h    0151A433    ;    //    slt x8 x3 x21      ====        slt s0, gp, s5
                                                  30'd    1491    : data = 32'h    27608A13    ;    //    addi x20 x1 630      ====        addi s4, ra, 630
                                                  30'd    1492    : data = 32'h    01B7D933    ;    //    srl x18 x15 x27      ====        srl s2, a5, s11
                                                  30'd    1493    : data = 32'h    E9F1C613    ;    //    xori x12 x3 -353      ====        xori a2, gp, -353
                                                  30'd    1494    : data = 32'h    013C8633    ;    //    add x12 x25 x19      ====        add a2, s9, s3
                                                  30'd    1495    : data = 32'h    415C8E33    ;    //    sub x28 x25 x21      ====        sub t3, s9, s5
                                                  30'd    1496    : data = 32'h    01073633    ;    //    sltu x12 x14 x16      ====        sltu a2, a4, a6
                                                  30'd    1497    : data = 32'h    3C7E4413    ;    //    xori x8 x28 967      ====        xori s0, t3, 967
                                                  30'd    1498    : data = 32'h    406489B3    ;    //    sub x19 x9 x6      ====        sub s3, s1, t1
                                                  30'd    1499    : data = 32'h    EC6BE013    ;    //    ori x0 x23 -314      ====        ori zero, s7, -314
                                                  30'd    1500    : data = 32'h    ABC56793    ;    //    ori x15 x10 -1348      ====        ori a5, a0, -1348
                                                  30'd    1501    : data = 32'h    7558FD93    ;    //    andi x27 x17 1877      ====        andi s11, a7, 1877
                                                  30'd    1502    : data = 32'h    A6CAB613    ;    //    sltiu x12 x21 -1428      ====        sltiu a2, s5, -1428
                                                  30'd    1503    : data = 32'h    413B5933    ;    //    sra x18 x22 x19      ====        sra s2, s6, s3
                                                  30'd    1504    : data = 32'h    40AF5D13    ;    //    srai x26 x30 10      ====        srai s10, t5, 10
                                                  30'd    1505    : data = 32'h    01A1C9B3    ;    //    xor x19 x3 x26      ====        xor s3, gp, s10
                                                  30'd    1506    : data = 32'h    B3C1E693    ;    //    ori x13 x3 -1220      ====        ori a3, gp, -1220
                                                  30'd    1507    : data = 32'h    00AFB4B3    ;    //    sltu x9 x31 x10      ====        sltu s1, t6, a0
                                                  30'd    1508    : data = 32'h    00D31EB3    ;    //    sll x29 x6 x13      ====        sll t4, t1, a3
                                                  30'd    1509    : data = 32'h    01B7CB33    ;    //    xor x22 x15 x27      ====        xor s6, a5, s11
                                                  30'd    1510    : data = 32'h    40630033    ;    //    sub x0 x6 x6      ====        sub zero, t1, t1
                                                  30'd    1511    : data = 32'h    01F8AD33    ;    //    slt x26 x17 x31      ====        slt s10, a7, t6
                                                  30'd    1512    : data = 32'h    00424333    ;    //    xor x6 x4 x4      ====        xor t1, tp, tp
                                                  30'd    1513    : data = 32'h    0057A3B3    ;    //    slt x7 x15 x5      ====        slt t2, a5, t0
                                                  30'd    1514    : data = 32'h    410450B3    ;    //    sra x1 x8 x16      ====        sra ra, s0, a6
                                                  30'd    1515    : data = 32'h    01705733    ;    //    srl x14 x0 x23      ====        srl a4, zero, s7
                                                  30'd    1516    : data = 32'h    011CDC93    ;    //    srli x25 x25 17      ====        srli s9, s9, 17
                                                  30'd    1517    : data = 32'h    83ECF393    ;    //    andi x7 x25 -1986      ====        andi t2, s9, -1986
                                                  30'd    1518    : data = 32'h    E93FBF93    ;    //    sltiu x31 x31 -365      ====        sltiu t6, t6, -365
                                                  30'd    1519    : data = 32'h    10B62293    ;    //    slti x5 x12 267      ====        slti t0, a2, 267
                                                  30'd    1520    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1521    : data = 32'h    973D4093    ;    //    xori x1 x26 -1677      ====        xori ra, s10, -1677
                                                  30'd    1522    : data = 32'h    ED454813    ;    //    xori x16 x10 -300      ====        xori a6, a0, -300
                                                  30'd    1523    : data = 32'h    DBEA3313    ;    //    sltiu x6 x20 -578      ====        sltiu t1, s4, -578
                                                  30'd    1524    : data = 32'h    0984ED13    ;    //    ori x26 x9 152      ====        ori s10, s1, 152
                                                  30'd    1525    : data = 32'h    01028FB3    ;    //    add x31 x5 x16      ====        add t6, t0, a6
                                                  30'd    1526    : data = 32'h    0139EAB3    ;    //    or x21 x19 x19      ====        or s5, s3, s3
                                                  30'd    1527    : data = 32'h    01CEACB3    ;    //    slt x25 x29 x28      ====        slt s9, t4, t3
                                                  30'd    1528    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1529    : data = 32'h    FBBE0E13    ;    //    addi x28 x28 -69      ====        addi t3, t3, -69
                                                  30'd    1530    : data = 32'h    016F5FB3    ;    //    srl x31 x30 x22      ====        srl t6, t5, s6
                                                  30'd    1531    : data = 32'h    404E5133    ;    //    sra x2 x28 x4      ====        sra sp, t3, tp
                                                  30'd    1532    : data = 32'h    014B9133    ;    //    sll x2 x23 x20      ====        sll sp, s7, s4
                                                  30'd    1533    : data = 32'h    000E2B33    ;    //    slt x22 x28 x0      ====        slt s6, t3, zero
                                                  30'd    1534    : data = 32'h    00A85E33    ;    //    srl x28 x16 x10      ====        srl t3, a6, a0
                                                  30'd    1535    : data = 32'h    A2883313    ;    //    sltiu x6 x16 -1496      ====        sltiu t1, a6, -1496
                                                  30'd    1536    : data = 32'h    403EDA93    ;    //    srai x21 x29 3      ====        srai s5, t4, 3
                                                  30'd    1537    : data = 32'h    004E59B3    ;    //    srl x19 x28 x4      ====        srl s3, t3, tp
                                                  30'd    1538    : data = 32'h    0002F933    ;    //    and x18 x5 x0      ====        and s2, t0, zero
                                                  30'd    1539    : data = 32'h    01A19733    ;    //    sll x14 x3 x26      ====        sll a4, gp, s10
                                                  30'd    1540    : data = 32'h    40070433    ;    //    sub x8 x14 x0      ====        sub s0, a4, zero
                                                  30'd    1541    : data = 32'h    002905B3    ;    //    add x11 x18 x2      ====        add a1, s2, sp
                                                  30'd    1542    : data = 32'h    0D5E4117    ;    //    auipc x2 54756      ====        auipc sp, 54756
                                                  30'd    1543    : data = 32'h    00280CB3    ;    //    add x25 x16 x2      ====        add s9, a6, sp
                                                  30'd    1544    : data = 32'h    017BCAB3    ;    //    xor x21 x23 x23      ====        xor s5, s7, s7
                                                  30'd    1545    : data = 32'h    0191BEB3    ;    //    sltu x29 x3 x25      ====        sltu t4, gp, s9
                                                  30'd    1546    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1547    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1548    : data = 32'h    41455793    ;    //    srai x15 x10 20      ====        srai a5, a0, 20
                                                  30'd    1549    : data = 32'h    01DD0133    ;    //    add x2 x26 x29      ====        add sp, s10, t4
                                                  30'd    1550    : data = 32'h    014D3733    ;    //    sltu x14 x26 x20      ====        sltu a4, s10, s4
                                                  30'd    1551    : data = 32'h    1A2D8793    ;    //    addi x15 x27 418      ====        addi a5, s11, 418
                                                  30'd    1552    : data = 32'h    1D4DE613    ;    //    ori x12 x27 468      ====        ori a2, s11, 468
                                                  30'd    1553    : data = 32'h    016384B3    ;    //    add x9 x7 x22      ====        add s1, t2, s6
                                                  30'd    1554    : data = 32'h    D3B70B93    ;    //    addi x23 x14 -709      ====        addi s7, a4, -709
                                                  30'd    1555    : data = 32'h    01BE1133    ;    //    sll x2 x28 x27      ====        sll sp, t3, s11
                                                  30'd    1556    : data = 32'h    01C11B13    ;    //    slli x22 x2 28      ====        slli s6, sp, 28
                                                  30'd    1557    : data = 32'h    ED883613    ;    //    sltiu x12 x16 -296      ====        sltiu a2, a6, -296
                                                  30'd    1558    : data = 32'h    B9943F93    ;    //    sltiu x31 x8 -1127      ====        sltiu t6, s0, -1127
                                                  30'd    1559    : data = 32'h    4520B093    ;    //    sltiu x1 x1 1106      ====        sltiu ra, ra, 1106
                                                  30'd    1560    : data = 32'h    00B2A733    ;    //    slt x14 x5 x11      ====        slt a4, t0, a1
                                                  30'd    1561    : data = 32'h    01DED693    ;    //    srli x13 x29 29      ====        srli a3, t4, 29
                                                  30'd    1562    : data = 32'h    F3493A93    ;    //    sltiu x21 x18 -204      ====        sltiu s5, s2, -204
                                                  30'd    1563    : data = 32'h    008335B3    ;    //    sltu x11 x6 x8      ====        sltu a1, t1, s0
                                                  30'd    1564    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1565    : data = 32'h    40435613    ;    //    srai x12 x6 4      ====        srai a2, t1, 4
                                                  30'd    1566    : data = 32'h    3884E813    ;    //    ori x16 x9 904      ====        ori a6, s1, 904
                                                  30'd    1567    : data = 32'h    50BB8593    ;    //    addi x11 x23 1291      ====        addi a1, s7, 1291
                                                  30'd    1568    : data = 32'h    01D0C433    ;    //    xor x8 x1 x29      ====        xor s0, ra, t4
                                                  30'd    1569    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1570    : data = 32'h    407209B3    ;    //    sub x19 x4 x7      ====        sub s3, tp, t2
                                                  30'd    1571    : data = 32'h    01ACA933    ;    //    slt x18 x25 x26      ====        slt s2, s9, s10
                                                  30'd    1572    : data = 32'h    0051B833    ;    //    sltu x16 x3 x5      ====        sltu a6, gp, t0
                                                  30'd    1573    : data = 32'h    0110C133    ;    //    xor x2 x1 x17      ====        xor sp, ra, a7
                                                  30'd    1574    : data = 32'h    41F8DE33    ;    //    sra x28 x17 x31      ====        sra t3, a7, t6
                                                  30'd    1575    : data = 32'h    00F305B3    ;    //    add x11 x6 x15      ====        add a1, t1, a5
                                                  30'd    1576    : data = 32'h    99AD0613    ;    //    addi x12 x26 -1638      ====        addi a2, s10, -1638
                                                  30'd    1577    : data = 32'h    00E4CD33    ;    //    xor x26 x9 x14      ====        xor s10, s1, a4
                                                  30'd    1578    : data = 32'h    01105C13    ;    //    srli x24 x0 17      ====        srli s8, zero, 17
                                                  30'd    1579    : data = 32'h    00125CB3    ;    //    srl x25 x4 x1      ====        srl s9, tp, ra
                                                  30'd    1580    : data = 32'h    61DE0B93    ;    //    addi x23 x28 1565      ====        addi s7, t3, 1565
                                                  30'd    1581    : data = 32'h    0FF82417    ;    //    auipc x8 65410      ====        auipc s0, 65410
                                                  30'd    1582    : data = 32'h    405903B3    ;    //    sub x7 x18 x5      ====        sub t2, s2, t0
                                                  30'd    1583    : data = 32'h    01D8AD33    ;    //    slt x26 x17 x29      ====        slt s10, a7, t4
                                                  30'd    1584    : data = 32'h    018ADBB3    ;    //    srl x23 x21 x24      ====        srl s7, s5, s8
                                                  30'd    1585    : data = 32'h    0196E133    ;    //    or x2 x13 x25      ====        or sp, a3, s9
                                                  30'd    1586    : data = 32'h    9198C613    ;    //    xori x12 x17 -1767      ====        xori a2, a7, -1767
                                                  30'd    1587    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1588    : data = 32'h    40848BB3    ;    //    sub x23 x9 x8      ====        sub s7, s1, s0
                                                  30'd    1589    : data = 32'h    007F6D33    ;    //    or x26 x30 x7      ====        or s10, t5, t2
                                                  30'd    1590    : data = 32'h    615CA113    ;    //    slti x2 x25 1557      ====        slti sp, s9, 1557
                                                  30'd    1591    : data = 32'h    00E10833    ;    //    add x16 x2 x14      ====        add a6, sp, a4
                                                  30'd    1592    : data = 32'h    00B5BC33    ;    //    sltu x24 x11 x11      ====        sltu s8, a1, a1
                                                  30'd    1593    : data = 32'h    01295D13    ;    //    srli x26 x18 18      ====        srli s10, s2, 18
                                                  30'd    1594    : data = 32'h    729A7493    ;    //    andi x9 x20 1833      ====        andi s1, s4, 1833
                                                  30'd    1595    : data = 32'h    B149CC13    ;    //    xori x24 x19 -1260      ====        xori s8, s3, -1260
                                                  30'd    1596    : data = 32'h    A5BC3917    ;    //    auipc x18 678851      ====        auipc s2, 678851
                                                  30'd    1597    : data = 32'h    0157D833    ;    //    srl x16 x15 x21      ====        srl a6, a5, s5
                                                  30'd    1598    : data = 32'h    4537ED37    ;    //    lui x26 283518      ====        lui s10, 283518
                                                  30'd    1599    : data = 32'h    70C87D93    ;    //    andi x27 x16 1804      ====        andi s11, a6, 1804
                                                  30'd    1600    : data = 32'h    01A11E13    ;    //    slli x28 x2 26      ====        slli t3, sp, 26
                                                  30'd    1601    : data = 32'h    ACF40093    ;    //    addi x1 x8 -1329      ====        addi ra, s0, -1329
                                                  30'd    1602    : data = 32'h    0045DB93    ;    //    srli x23 x11 4      ====        srli s7, a1, 4
                                                  30'd    1603    : data = 32'h    403AD733    ;    //    sra x14 x21 x3      ====        sra a4, s5, gp
                                                  30'd    1604    : data = 32'h    019B5C33    ;    //    srl x24 x22 x25      ====        srl s8, s6, s9
                                                  30'd    1605    : data = 32'h    A38B8613    ;    //    addi x12 x23 -1480      ====        addi a2, s7, -1480
                                                  30'd    1606    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1607    : data = 32'h    32020E13    ;    //    addi x28 x4 800      ====        addi t3, tp, 800
                                                  30'd    1608    : data = 32'h    00975EB3    ;    //    srl x29 x14 x9      ====        srl t4, a4, s1
                                                  30'd    1609    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1610    : data = 32'h    01730A33    ;    //    add x20 x6 x23      ====        add s4, t1, s7
                                                  30'd    1611    : data = 32'h    9165AD93    ;    //    slti x27 x11 -1770      ====        slti s11, a1, -1770
                                                  30'd    1612    : data = 32'h    82C60913    ;    //    addi x18 x12 -2004      ====        addi s2, a2, -2004
                                                  30'd    1613    : data = 32'h    0DBA2A93    ;    //    slti x21 x20 219      ====        slti s5, s4, 219
                                                  30'd    1614    : data = 32'h    01A7B1B3    ;    //    sltu x3 x15 x26      ====        sltu gp, a5, s10
                                                  30'd    1615    : data = 32'h    856B2093    ;    //    slti x1 x22 -1962      ====        slti ra, s6, -1962
                                                  30'd    1616    : data = 32'h    4009D133    ;    //    sra x2 x19 x0      ====        sra sp, s3, zero
                                                  30'd    1617    : data = 32'h    40925133    ;    //    sra x2 x4 x9      ====        sra sp, tp, s1
                                                  30'd    1618    : data = 32'h    00EBD913    ;    //    srli x18 x23 14      ====        srli s2, s7, 14
                                                  30'd    1619    : data = 32'h    00779C93    ;    //    slli x25 x15 7      ====        slli s9, a5, 7
                                                  30'd    1620    : data = 32'h    706B8713    ;    //    addi x14 x23 1798      ====        addi a4, s7, 1798
                                                  30'd    1621    : data = 32'h    EA016893    ;    //    ori x17 x2 -352      ====        ori a7, sp, -352
                                                  30'd    1622    : data = 32'h    01036AB3    ;    //    or x21 x6 x16      ====        or s5, t1, a6
                                                  30'd    1623    : data = 32'h    48B1F893    ;    //    andi x17 x3 1163      ====        andi a7, gp, 1163
                                                  30'd    1624    : data = 32'h    01D1D433    ;    //    srl x8 x3 x29      ====        srl s0, gp, t4
                                                  30'd    1625    : data = 32'h    40CED993    ;    //    srai x19 x29 12      ====        srai s3, t4, 12
                                                  30'd    1626    : data = 32'h    0005D613    ;    //    srli x12 x11 0      ====        srli a2, a1, 0
                                                  30'd    1627    : data = 32'h    00D59293    ;    //    slli x5 x11 13      ====        slli t0, a1, 13
                                                  30'd    1628    : data = 32'h    40FBD6B3    ;    //    sra x13 x23 x15      ====        sra a3, s7, a5
                                                  30'd    1629    : data = 32'h    91717293    ;    //    andi x5 x2 -1769      ====        andi t0, sp, -1769
                                                  30'd    1630    : data = 32'h    01342B33    ;    //    slt x22 x8 x19      ====        slt s6, s0, s3
                                                  30'd    1631    : data = 32'h    01479013    ;    //    slli x0 x15 20      ====        slli zero, a5, 20
                                                  30'd    1632    : data = 32'h    01E8DCB3    ;    //    srl x25 x17 x30      ====        srl s9, a7, t5
                                                  30'd    1633    : data = 32'h    01F3B133    ;    //    sltu x2 x7 x31      ====        sltu sp, t2, t6
                                                  30'd    1634    : data = 32'h    46217293    ;    //    andi x5 x2 1122      ====        andi t0, sp, 1122
                                                  30'd    1635    : data = 32'h    01F9E2B3    ;    //    or x5 x19 x31      ====        or t0, s3, t6
                                                  30'd    1636    : data = 32'h    0157B6B3    ;    //    sltu x13 x15 x21      ====        sltu a3, a5, s5
                                                  30'd    1637    : data = 32'h    420A0997    ;    //    auipc x19 270496      ====        auipc s3, 270496
                                                  30'd    1638    : data = 32'h    B55FCD13    ;    //    xori x26 x31 -1195      ====        xori s10, t6, -1195
                                                  30'd    1639    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1640    : data = 32'h    408F5793    ;    //    srai x15 x30 8      ====        srai a5, t5, 8
                                                  30'd    1641    : data = 32'h    2A88A293    ;    //    slti x5 x17 680      ====        slti t0, a7, 680
                                                  30'd    1642    : data = 32'h    FD65C613    ;    //    xori x12 x11 -42      ====        xori a2, a1, -42
                                                  30'd    1643    : data = 32'h    B7A14997    ;    //    auipc x19 752148      ====        auipc s3, 752148
                                                  30'd    1644    : data = 32'h    F2C333B7    ;    //    lui x7 994355      ====        lui t2, 994355
                                                  30'd    1645    : data = 32'h    00824833    ;    //    xor x16 x4 x8      ====        xor a6, tp, s0
                                                  30'd    1646    : data = 32'h    01BECEB3    ;    //    xor x29 x29 x27      ====        xor t4, t4, s11
                                                  30'd    1647    : data = 32'h    00BF9293    ;    //    slli x5 x31 11      ====        slli t0, t6, 11
                                                  30'd    1648    : data = 32'h    00DE45B3    ;    //    xor x11 x28 x13      ====        xor a1, t3, a3
                                                  30'd    1649    : data = 32'h    410E5DB3    ;    //    sra x27 x28 x16      ====        sra s11, t3, a6
                                                  30'd    1650    : data = 32'h    00D34FB3    ;    //    xor x31 x6 x13      ====        xor t6, t1, a3
                                                  30'd    1651    : data = 32'h    01470BB3    ;    //    add x23 x14 x20      ====        add s7, a4, s4
                                                  30'd    1652    : data = 32'h    0914C893    ;    //    xori x17 x9 145      ====        xori a7, s1, 145
                                                  30'd    1653    : data = 32'h    191ABB93    ;    //    sltiu x23 x21 401      ====        sltiu s7, s5, 401
                                                  30'd    1654    : data = 32'h    01C3EEB3    ;    //    or x29 x7 x28      ====        or t4, t2, t3
                                                  30'd    1655    : data = 32'h    AFCAFF93    ;    //    andi x31 x21 -1284      ====        andi t6, s5, -1284
                                                  30'd    1656    : data = 32'h    017C69B3    ;    //    or x19 x24 x23      ====        or s3, s8, s7
                                                  30'd    1657    : data = 32'h    00233D33    ;    //    sltu x26 x6 x2      ====        sltu s10, t1, sp
                                                  30'd    1658    : data = 32'h    0155A5B3    ;    //    slt x11 x11 x21      ====        slt a1, a1, s5
                                                  30'd    1659    : data = 32'h    00794C33    ;    //    xor x24 x18 x7      ====        xor s8, s2, t2
                                                  30'd    1660    : data = 32'h    0047C933    ;    //    xor x18 x15 x4      ====        xor s2, a5, tp
                                                  30'd    1661    : data = 32'h    40BDDA93    ;    //    srai x21 x27 11      ====        srai s5, s11, 11
                                                  30'd    1662    : data = 32'h    52B17D13    ;    //    andi x26 x2 1323      ====        andi s10, sp, 1323
                                                  30'd    1663    : data = 32'h    402684B3    ;    //    sub x9 x13 x2      ====        sub s1, a3, sp
                                                  30'd    1664    : data = 32'h    01344733    ;    //    xor x14 x8 x19      ====        xor a4, s0, s3
                                                  30'd    1665    : data = 32'h    00C75E33    ;    //    srl x28 x14 x12      ====        srl t3, a4, a2
                                                  30'd    1666    : data = 32'h    01E4D733    ;    //    srl x14 x9 x30      ====        srl a4, s1, t5
                                                  30'd    1667    : data = 32'h    01557433    ;    //    and x8 x10 x21      ====        and s0, a0, s5
                                                  30'd    1668    : data = 32'h    ADA3E493    ;    //    ori x9 x7 -1318      ====        ori s1, t2, -1318
                                                  30'd    1669    : data = 32'h    413C5F93    ;    //    srai x31 x24 19      ====        srai t6, s8, 19
                                                  30'd    1670    : data = 32'h    01B479B3    ;    //    and x19 x8 x27      ====        and s3, s0, s11
                                                  30'd    1671    : data = 32'h    001B5833    ;    //    srl x16 x22 x1      ====        srl a6, s6, ra
                                                  30'd    1672    : data = 32'h    01F1A9B3    ;    //    slt x19 x3 x31      ====        slt s3, gp, t6
                                                  30'd    1673    : data = 32'h    770B6D37    ;    //    lui x26 487606      ====        lui s10, 487606
                                                  30'd    1674    : data = 32'h    08B6FC93    ;    //    andi x25 x13 139      ====        andi s9, a3, 139
                                                  30'd    1675    : data = 32'h    793E3A13    ;    //    sltiu x20 x28 1939      ====        sltiu s4, t3, 1939
                                                  30'd    1676    : data = 32'h    01FB06B3    ;    //    add x13 x22 x31      ====        add a3, s6, t6
                                                  30'd    1677    : data = 32'h    01FA9E33    ;    //    sll x28 x21 x31      ====        sll t3, s5, t6
                                                  30'd    1678    : data = 32'h    45CE8013    ;    //    addi x0 x29 1116      ====        addi zero, t4, 1116
                                                  30'd    1679    : data = 32'h    B89DAC93    ;    //    slti x25 x27 -1143      ====        slti s9, s11, -1143
                                                  30'd    1680    : data = 32'h    0141FFB3    ;    //    and x31 x3 x20      ====        and t6, gp, s4
                                                  30'd    1681    : data = 32'h    F66F7013    ;    //    andi x0 x30 -154      ====        andi zero, t5, -154
                                                  30'd    1682    : data = 32'h    01251793    ;    //    slli x15 x10 18      ====        slli a5, a0, 18
                                                  30'd    1683    : data = 32'h    DDCFF8B7    ;    //    lui x17 908543      ====        lui a7, 908543
                                                  30'd    1684    : data = 32'h    0B4D7737    ;    //    lui x14 46295      ====        lui a4, 46295
                                                  30'd    1685    : data = 32'h    01722033    ;    //    slt x0 x4 x23      ====        slt zero, tp, s7
                                                  30'd    1686    : data = 32'h    01375693    ;    //    srli x13 x14 19      ====        srli a3, a4, 19
                                                  30'd    1687    : data = 32'h    00810B33    ;    //    add x22 x2 x8      ====        add s6, sp, s0
                                                  30'd    1688    : data = 32'h    013A8733    ;    //    add x14 x21 x19      ====        add a4, s5, s3
                                                  30'd    1689    : data = 32'h    41078C33    ;    //    sub x24 x15 x16      ====        sub s8, a5, a6
                                                  30'd    1690    : data = 32'h    AEAAD817    ;    //    auipc x16 715437      ====        auipc a6, 715437
                                                  30'd    1691    : data = 32'h    00FF5713    ;    //    srli x14 x30 15      ====        srli a4, t5, 15
                                                  30'd    1692    : data = 32'h    01975AB3    ;    //    srl x21 x14 x25      ====        srl s5, a4, s9
                                                  30'd    1693    : data = 32'h    0048EAB3    ;    //    or x21 x17 x4      ====        or s5, a7, tp
                                                  30'd    1694    : data = 32'h    0809FE17    ;    //    auipc x28 32927      ====        auipc t3, 32927
                                                  30'd    1695    : data = 32'h    40A9DFB3    ;    //    sra x31 x19 x10      ====        sra t6, s3, a0
                                                  30'd    1696    : data = 32'h    01411C93    ;    //    slli x25 x2 20      ====        slli s9, sp, 20
                                                  30'd    1697    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1698    : data = 32'h    00CB86B3    ;    //    add x13 x23 x12      ====        add a3, s7, a2
                                                  30'd    1699    : data = 32'h    BCAE4293    ;    //    xori x5 x28 -1078      ====        xori t0, t3, -1078
                                                  30'd    1700    : data = 32'h    AE1AAD13    ;    //    slti x26 x21 -1311      ====        slti s10, s5, -1311
                                                  30'd    1701    : data = 32'h    B5A04DB7    ;    //    lui x27 743940      ====        lui s11, 743940
                                                  30'd    1702    : data = 32'h    8666FE93    ;    //    andi x29 x13 -1946      ====        andi t4, a3, -1946
                                                  30'd    1703    : data = 32'h    0095C9B3    ;    //    xor x19 x11 x9      ====        xor s3, a1, s1
                                                  30'd    1704    : data = 32'h    4017D813    ;    //    srai x16 x15 1      ====        srai a6, a5, 1
                                                  30'd    1705    : data = 32'h    41FC0633    ;    //    sub x12 x24 x31      ====        sub a2, s8, t6
                                                  30'd    1706    : data = 32'h    0191DD33    ;    //    srl x26 x3 x25      ====        srl s10, gp, s9
                                                  30'd    1707    : data = 32'h    01EE71B3    ;    //    and x3 x28 x30      ====        and gp, t3, t5
                                                  30'd    1708    : data = 32'h    7123AE13    ;    //    slti x28 x7 1810      ====        slti t3, t2, 1810
                                                  30'd    1709    : data = 32'h    04DC7613    ;    //    andi x12 x24 77      ====        andi a2, s8, 77
                                                  30'd    1710    : data = 32'h    B4A88D93    ;    //    addi x27 x17 -1206      ====        addi s11, a7, -1206
                                                  30'd    1711    : data = 32'h    0049D633    ;    //    srl x12 x19 x4      ====        srl a2, s3, tp
                                                  30'd    1712    : data = 32'h    016B1D13    ;    //    slli x26 x22 22      ====        slli s10, s6, 22
                                                  30'd    1713    : data = 32'h    00F39013    ;    //    slli x0 x7 15      ====        slli zero, t2, 15
                                                  30'd    1714    : data = 32'h    41818033    ;    //    sub x0 x3 x24      ====        sub zero, gp, s8
                                                  30'd    1715    : data = 32'h    01BEF7B3    ;    //    and x15 x29 x27      ====        and a5, t4, s11
                                                  30'd    1716    : data = 32'h    EEBB2337    ;    //    lui x6 977842      ====        lui t1, 977842
                                                  30'd    1717    : data = 32'h    011D2BB3    ;    //    slt x23 x26 x17      ====        slt s7, s10, a7
                                                  30'd    1718    : data = 32'h    F6D73813    ;    //    sltiu x16 x14 -147      ====        sltiu a6, a4, -147
                                                  30'd    1719    : data = 32'h    01E2D693    ;    //    srli x13 x5 30      ====        srli a3, t0, 30
                                                  30'd    1720    : data = 32'h    015B7833    ;    //    and x16 x22 x21      ====        and a6, s6, s5
                                                  30'd    1721    : data = 32'h    0100CFB3    ;    //    xor x31 x1 x16      ====        xor t6, ra, a6
                                                  30'd    1722    : data = 32'h    F94B7113    ;    //    andi x2 x22 -108      ====        andi sp, s6, -108
                                                  30'd    1723    : data = 32'h    00D2FEB3    ;    //    and x29 x5 x13      ====        and t4, t0, a3
                                                  30'd    1724    : data = 32'h    0099D113    ;    //    srli x2 x19 9      ====        srli sp, s3, 9
                                                  30'd    1725    : data = 32'h    01C2BCB3    ;    //    sltu x25 x5 x28      ====        sltu s9, t0, t3
                                                  30'd    1726    : data = 32'h    173695B7    ;    //    lui x11 95081      ====        lui a1, 95081
                                                  30'd    1727    : data = 32'h    49D40437    ;    //    lui x8 302400      ====        lui s0, 302400
                                                  30'd    1728    : data = 32'h    0070B0B3    ;    //    sltu x1 x1 x7      ====        sltu ra, ra, t2
                                                  30'd    1729    : data = 32'h    00211A13    ;    //    slli x20 x2 2      ====        slli s4, sp, 2
                                                  30'd    1730    : data = 32'h    3EE9AF93    ;    //    slti x31 x19 1006      ====        slti t6, s3, 1006
                                                  30'd    1731    : data = 32'h    01B6ACB3    ;    //    slt x25 x13 x27      ====        slt s9, a3, s11
                                                  30'd    1732    : data = 32'h    014A78B3    ;    //    and x17 x20 x20      ====        and a7, s4, s4
                                                  30'd    1733    : data = 32'h    015DDEB3    ;    //    srl x29 x27 x21      ====        srl t4, s11, s5
                                                  30'd    1734    : data = 32'h    009DEFB3    ;    //    or x31 x27 x9      ====        or t6, s11, s1
                                                  30'd    1735    : data = 32'h    40B1D2B3    ;    //    sra x5 x3 x11      ====        sra t0, gp, a1
                                                  30'd    1736    : data = 32'h    4C297713    ;    //    andi x14 x18 1218      ====        andi a4, s2, 1218
                                                  30'd    1737    : data = 32'h    8DAD5FB7    ;    //    lui x31 580309      ====        lui t6, 580309
                                                  30'd    1738    : data = 32'h    012AA433    ;    //    slt x8 x21 x18      ====        slt s0, s5, s2
                                                  30'd    1739    : data = 32'h    0139EC33    ;    //    or x24 x19 x19      ====        or s8, s3, s3
                                                  30'd    1740    : data = 32'h    BA357913    ;    //    andi x18 x10 -1117      ====        andi s2, a0, -1117
                                                  30'd    1741    : data = 32'h    010319B3    ;    //    sll x19 x6 x16      ====        sll s3, t1, a6
                                                  30'd    1742    : data = 32'h    40328733    ;    //    sub x14 x5 x3      ====        sub a4, t0, gp
                                                  30'd    1743    : data = 32'h    CF1E0D13    ;    //    addi x26 x28 -783      ====        addi s10, t3, -783
                                                  30'd    1744    : data = 32'h    769BA813    ;    //    slti x16 x23 1897      ====        slti a6, s7, 1897
                                                  30'd    1745    : data = 32'h    00BE8C33    ;    //    add x24 x29 x11      ====        add s8, t4, a1
                                                  30'd    1746    : data = 32'h    017A5B33    ;    //    srl x22 x20 x23      ====        srl s6, s4, s7
                                                  30'd    1747    : data = 32'h    0075A133    ;    //    slt x2 x11 x7      ====        slt sp, a1, t2
                                                  30'd    1748    : data = 32'h    CEA0CE13    ;    //    xori x28 x1 -790      ====        xori t3, ra, -790
                                                  30'd    1749    : data = 32'h    5D8F3813    ;    //    sltiu x16 x30 1496      ====        sltiu a6, t5, 1496
                                                  30'd    1750    : data = 32'h    5328CB93    ;    //    xori x23 x17 1330      ====        xori s7, a7, 1330
                                                  30'd    1751    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1752    : data = 32'h    009EB833    ;    //    sltu x16 x29 x9      ====        sltu a6, t4, s1
                                                  30'd    1753    : data = 32'h    00F14433    ;    //    xor x8 x2 x15      ====        xor s0, sp, a5
                                                  30'd    1754    : data = 32'h    D5944D13    ;    //    xori x26 x8 -679      ====        xori s10, s0, -679
                                                  30'd    1755    : data = 32'h    004CB5B3    ;    //    sltu x11 x25 x4      ====        sltu a1, s9, tp
                                                  30'd    1756    : data = 32'h    DD264293    ;    //    xori x5 x12 -558      ====        xori t0, a2, -558
                                                  30'd    1757    : data = 32'h    05827113    ;    //    andi x2 x4 88      ====        andi sp, tp, 88
                                                  30'd    1758    : data = 32'h    69E25E97    ;    //    auipc x29 433701      ====        auipc t4, 433701
                                                  30'd    1759    : data = 32'h    016BAFB3    ;    //    slt x31 x23 x22      ====        slt t6, s7, s6
                                                  30'd    1760    : data = 32'h    A7508393    ;    //    addi x7 x1 -1419      ====        addi t2, ra, -1419
                                                  30'd    1761    : data = 32'h    C3030793    ;    //    addi x15 x6 -976      ====        addi a5, t1, -976
                                                  30'd    1762    : data = 32'h    01537033    ;    //    and x0 x6 x21      ====        and zero, t1, s5
                                                  30'd    1763    : data = 32'h    23C10393    ;    //    addi x7 x2 572      ====        addi t2, sp, 572
                                                  30'd    1764    : data = 32'h    0136DB93    ;    //    srli x23 x13 19      ====        srli s7, a3, 19
                                                  30'd    1765    : data = 32'h    40925993    ;    //    srai x19 x4 9      ====        srai s3, tp, 9
                                                  30'd    1766    : data = 32'h    E77CCE13    ;    //    xori x28 x25 -393      ====        xori t3, s9, -393
                                                  30'd    1767    : data = 32'h    400AD633    ;    //    sra x12 x21 x0      ====        sra a2, s5, zero
                                                  30'd    1768    : data = 32'h    BACDE117    ;    //    auipc x2 765150      ====        auipc sp, 765150
                                                  30'd    1769    : data = 32'h    2537E013    ;    //    ori x0 x15 595      ====        ori zero, a5, 595
                                                  30'd    1770    : data = 32'h    01E29B93    ;    //    slli x23 x5 30      ====        slli s7, t0, 30
                                                  30'd    1771    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1772    : data = 32'h    25A02913    ;    //    slti x18 x0 602      ====        slti s2, zero, 602
                                                  30'd    1773    : data = 32'h    19BD3D93    ;    //    sltiu x27 x26 411      ====        sltiu s11, s10, 411
                                                  30'd    1774    : data = 32'h    00C35B13    ;    //    srli x22 x6 12      ====        srli s6, t1, 12
                                                  30'd    1775    : data = 32'h    0145DD33    ;    //    srl x26 x11 x20      ====        srl s10, a1, s4
                                                  30'd    1776    : data = 32'h    015ED813    ;    //    srli x16 x29 21      ====        srli a6, t4, 21
                                                  30'd    1777    : data = 32'h    01D04033    ;    //    xor x0 x0 x29      ====        xor zero, zero, t4
                                                  30'd    1778    : data = 32'h    00A29CB3    ;    //    sll x25 x5 x10      ====        sll s9, t0, a0
                                                  30'd    1779    : data = 32'h    015D03B3    ;    //    add x7 x26 x21      ====        add t2, s10, s5
                                                  30'd    1780    : data = 32'h    01E36933    ;    //    or x18 x6 x30      ====        or s2, t1, t5
                                                  30'd    1781    : data = 32'h    014E7933    ;    //    and x18 x28 x20      ====        and s2, t3, s4
                                                  30'd    1782    : data = 32'h    5A478C13    ;    //    addi x24 x15 1444      ====        addi s8, a5, 1444
                                                  30'd    1783    : data = 32'h    EB1C3A93    ;    //    sltiu x21 x24 -335      ====        sltiu s5, s8, -335
                                                  30'd    1784    : data = 32'h    0060F033    ;    //    and x0 x1 x6      ====        and zero, ra, t1
                                                  30'd    1785    : data = 32'h    01AC47B3    ;    //    xor x15 x24 x26      ====        xor a5, s8, s10
                                                  30'd    1786    : data = 32'h    40745393    ;    //    srai x7 x8 7      ====        srai t2, s0, 7
                                                  30'd    1787    : data = 32'h    01F94433    ;    //    xor x8 x18 x31      ====        xor s0, s2, t6
                                                  30'd    1788    : data = 32'h    0F92AB93    ;    //    slti x23 x5 249      ====        slti s7, t0, 249
                                                  30'd    1789    : data = 32'h    00F12E33    ;    //    slt x28 x2 x15      ====        slt t3, sp, a5
                                                  30'd    1790    : data = 32'h    002AA5B3    ;    //    slt x11 x21 x2      ====        slt a1, s5, sp
                                                  30'd    1791    : data = 32'h    01D627B3    ;    //    slt x15 x12 x29      ====        slt a5, a2, t4
                                                  30'd    1792    : data = 32'h    C37C1017    ;    //    auipc x0 800705      ====        auipc zero, 800705
                                                  30'd    1793    : data = 32'h    01AEBEB3    ;    //    sltu x29 x29 x26      ====        sltu t4, t4, s10
                                                  30'd    1794    : data = 32'h    013E0833    ;    //    add x16 x28 x19      ====        add a6, t3, s3
                                                  30'd    1795    : data = 32'h    8F9D8013    ;    //    addi x0 x27 -1799      ====        addi zero, s11, -1799
                                                  30'd    1796    : data = 32'h    26AE6D13    ;    //    ori x26 x28 618      ====        ori s10, t3, 618
                                                  30'd    1797    : data = 32'h    009F9B13    ;    //    slli x22 x31 9      ====        slli s6, t6, 9
                                                  30'd    1798    : data = 32'h    00FB6433    ;    //    or x8 x22 x15      ====        or s0, s6, a5
                                                  30'd    1799    : data = 32'h    01907CB3    ;    //    and x25 x0 x25      ====        and s9, zero, s9
                                                  30'd    1800    : data = 32'h    6148F313    ;    //    andi x6 x17 1556      ====        andi t1, a7, 1556
                                                  30'd    1801    : data = 32'h    407B0033    ;    //    sub x0 x22 x7      ====        sub zero, s6, t2
                                                  30'd    1802    : data = 32'h    01CB7033    ;    //    and x0 x22 x28      ====        and zero, s6, t3
                                                  30'd    1803    : data = 32'h    00A95BB3    ;    //    srl x23 x18 x10      ====        srl s7, s2, a0
                                                  30'd    1804    : data = 32'h    E8268A37    ;    //    lui x20 950888      ====        lui s4, 950888
                                                  30'd    1805    : data = 32'h    415D0C33    ;    //    sub x24 x26 x21      ====        sub s8, s10, s5
                                                  30'd    1806    : data = 32'h    4006DC93    ;    //    srai x25 x13 0      ====        srai s9, a3, 0
                                                  30'd    1807    : data = 32'h    017A1793    ;    //    slli x15 x20 23      ====        slli a5, s4, 23
                                                  30'd    1808    : data = 32'h    B54A4093    ;    //    xori x1 x20 -1196      ====        xori ra, s4, -1196
                                                  30'd    1809    : data = 32'h    411BD193    ;    //    srai x3 x23 17      ====        srai gp, s7, 17
                                                  30'd    1810    : data = 32'h    01349333    ;    //    sll x6 x9 x19      ====        sll t1, s1, s3
                                                  30'd    1811    : data = 32'h    011DC433    ;    //    xor x8 x27 x17      ====        xor s0, s11, a7
                                                  30'd    1812    : data = 32'h    0161E0B3    ;    //    or x1 x3 x22      ====        or ra, gp, s6
                                                  30'd    1813    : data = 32'h    77617717    ;    //    auipc x14 488983      ====        auipc a4, 488983
                                                  30'd    1814    : data = 32'h    010DFE33    ;    //    and x28 x27 x16      ====        and t3, s11, a6
                                                  30'd    1815    : data = 32'h    0138DE93    ;    //    srli x29 x17 19      ====        srli t4, a7, 19
                                                  30'd    1816    : data = 32'h    C7F42893    ;    //    slti x17 x8 -897      ====        slti a7, s0, -897
                                                  30'd    1817    : data = 32'h    0102B9B3    ;    //    sltu x19 x5 x16      ====        sltu s3, t0, a6
                                                  30'd    1818    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1819    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1820    : data = 32'h    41525D13    ;    //    srai x26 x4 21      ====        srai s10, tp, 21
                                                  30'd    1821    : data = 32'h    307F0E97    ;    //    auipc x29 198640      ====        auipc t4, 198640
                                                  30'd    1822    : data = 32'h    00899113    ;    //    slli x2 x19 8      ====        slli sp, s3, 8
                                                  30'd    1823    : data = 32'h    3DCE6113    ;    //    ori x2 x28 988      ====        ori sp, t3, 988
                                                  30'd    1824    : data = 32'h    000A1133    ;    //    sll x2 x20 x0      ====        sll sp, s4, zero
                                                  30'd    1825    : data = 32'h    EBBFEB93    ;    //    ori x23 x31 -325      ====        ori s7, t6, -325
                                                  30'd    1826    : data = 32'h    0EACE013    ;    //    ori x0 x25 234      ====        ori zero, s9, 234
                                                  30'd    1827    : data = 32'h    786A3593    ;    //    sltiu x11 x20 1926      ====        sltiu a1, s4, 1926
                                                  30'd    1828    : data = 32'h    A9B52D93    ;    //    slti x27 x10 -1381      ====        slti s11, a0, -1381
                                                  30'd    1829    : data = 32'h    00F82CB3    ;    //    slt x25 x16 x15      ====        slt s9, a6, a5
                                                  30'd    1830    : data = 32'h    00EA2C33    ;    //    slt x24 x20 x14      ====        slt s8, s4, a4
                                                  30'd    1831    : data = 32'h    01225833    ;    //    srl x16 x4 x18      ====        srl a6, tp, s2
                                                  30'd    1832    : data = 32'h    E9677F93    ;    //    andi x31 x14 -362      ====        andi t6, a4, -362
                                                  30'd    1833    : data = 32'h    004C2B33    ;    //    slt x22 x24 x4      ====        slt s6, s8, tp
                                                  30'd    1834    : data = 32'h    00B9A6B3    ;    //    slt x13 x19 x11      ====        slt a3, s3, a1
                                                  30'd    1835    : data = 32'h    4093DC13    ;    //    srai x24 x7 9      ====        srai s8, t2, 9
                                                  30'd    1836    : data = 32'h    0C61A913    ;    //    slti x18 x3 198      ====        slti s2, gp, 198
                                                  30'd    1837    : data = 32'h    399FAD13    ;    //    slti x26 x31 921      ====        slti s10, t6, 921
                                                  30'd    1838    : data = 32'h    007F5893    ;    //    srli x17 x30 7      ====        srli a7, t5, 7
                                                  30'd    1839    : data = 32'h    B19DE413    ;    //    ori x8 x27 -1255      ====        ori s0, s11, -1255
                                                  30'd    1840    : data = 32'h    40A581B3    ;    //    sub x3 x11 x10      ====        sub gp, a1, a0
                                                  30'd    1841    : data = 32'h    00D7CDB3    ;    //    xor x27 x15 x13      ====        xor s11, a5, a3
                                                  30'd    1842    : data = 32'h    000345B3    ;    //    xor x11 x6 x0      ====        xor a1, t1, zero
                                                  30'd    1843    : data = 32'h    0076B933    ;    //    sltu x18 x13 x7      ====        sltu s2, a3, t2
                                                  30'd    1844    : data = 32'h    008BAD33    ;    //    slt x26 x23 x8      ====        slt s10, s7, s0
                                                  30'd    1845    : data = 32'h    005194B3    ;    //    sll x9 x3 x5      ====        sll s1, gp, t0
                                                  30'd    1846    : data = 32'h    010AD833    ;    //    srl x16 x21 x16      ====        srl a6, s5, a6
                                                  30'd    1847    : data = 32'h    411E5D93    ;    //    srai x27 x28 17      ====        srai s11, t3, 17
                                                  30'd    1848    : data = 32'h    4098D5B3    ;    //    sra x11 x17 x9      ====        sra a1, a7, s1
                                                  30'd    1849    : data = 32'h    00825D13    ;    //    srli x26 x4 8      ====        srli s10, tp, 8
                                                  30'd    1850    : data = 32'h    A98C0593    ;    //    addi x11 x24 -1384      ====        addi a1, s8, -1384
                                                  30'd    1851    : data = 32'h    01861293    ;    //    slli x5 x12 24      ====        slli t0, a2, 24
                                                  30'd    1852    : data = 32'h    984F0493    ;    //    addi x9 x30 -1660      ====        addi s1, t5, -1660
                                                  30'd    1853    : data = 32'h    BFF2AC13    ;    //    slti x24 x5 -1025      ====        slti s8, t0, -1025
                                                  30'd    1854    : data = 32'h    40DDD493    ;    //    srai x9 x27 13      ====        srai s1, s11, 13
                                                  30'd    1855    : data = 32'h    01776B33    ;    //    or x22 x14 x23      ====        or s6, a4, s7
                                                  30'd    1856    : data = 32'h    01981133    ;    //    sll x2 x16 x25      ====        sll sp, a6, s9
                                                  30'd    1857    : data = 32'h    4552A613    ;    //    slti x12 x5 1109      ====        slti a2, t0, 1109
                                                  30'd    1858    : data = 32'h    40C4D013    ;    //    srai x0 x9 12      ====        srai zero, s1, 12
                                                  30'd    1859    : data = 32'h    01D76033    ;    //    or x0 x14 x29      ====        or zero, a4, t4
                                                  30'd    1860    : data = 32'h    220C6493    ;    //    ori x9 x24 544      ====        ori s1, s8, 544
                                                  30'd    1861    : data = 32'h    1EA66C93    ;    //    ori x25 x12 490      ====        ori s9, a2, 490
                                                  30'd    1862    : data = 32'h    99F13E13    ;    //    sltiu x28 x2 -1633      ====        sltiu t3, sp, -1633
                                                  30'd    1863    : data = 32'h    01F442B3    ;    //    xor x5 x8 x31      ====        xor t0, s0, t6
                                                  30'd    1864    : data = 32'h    01FB96B3    ;    //    sll x13 x23 x31      ====        sll a3, s7, t6
                                                  30'd    1865    : data = 32'h    62417837    ;    //    lui x16 402455      ====        lui a6, 402455
                                                  30'd    1866    : data = 32'h    41CF89B3    ;    //    sub x19 x31 x28      ====        sub s3, t6, t3
                                                  30'd    1867    : data = 32'h    00F372B3    ;    //    and x5 x6 x15      ====        and t0, t1, a5
                                                  30'd    1868    : data = 32'h    405056B3    ;    //    sra x13 x0 x5      ====        sra a3, zero, t0
                                                  30'd    1869    : data = 32'h    2F81CC97    ;    //    auipc x25 194588      ====        auipc s9, 194588
                                                  30'd    1870    : data = 32'h    000E9293    ;    //    slli x5 x29 0      ====        slli t0, t4, 0
                                                  30'd    1871    : data = 32'h    00D3D933    ;    //    srl x18 x7 x13      ====        srl s2, t2, a3
                                                  30'd    1872    : data = 32'h    00571293    ;    //    slli x5 x14 5      ====        slli t0, a4, 5
                                                  30'd    1873    : data = 32'h    012EBD33    ;    //    sltu x26 x29 x18      ====        sltu s10, t4, s2
                                                  30'd    1874    : data = 32'h    4019D6B3    ;    //    sra x13 x19 x1      ====        sra a3, s3, ra
                                                  30'd    1875    : data = 32'h    00079A33    ;    //    sll x20 x15 x0      ====        sll s4, a5, zero
                                                  30'd    1876    : data = 32'h    404A5593    ;    //    srai x11 x20 4      ====        srai a1, s4, 4
                                                  30'd    1877    : data = 32'h    0023CBB3    ;    //    xor x23 x7 x2      ====        xor s7, t2, sp
                                                  30'd    1878    : data = 32'h    001CD713    ;    //    srli x14 x25 1      ====        srli a4, s9, 1
                                                  30'd    1879    : data = 32'h    00C9AD33    ;    //    slt x26 x19 x12      ====        slt s10, s3, a2
                                                  30'd    1880    : data = 32'h    75AEB813    ;    //    sltiu x16 x29 1882      ====        sltiu a6, t4, 1882
                                                  30'd    1881    : data = 32'h    D4C10493    ;    //    addi x9 x2 -692      ====        addi s1, sp, -692
                                                  30'd    1882    : data = 32'h    6FC06293    ;    //    ori x5 x0 1788      ====        ori t0, zero, 1788
                                                  30'd    1883    : data = 32'h    016592B3    ;    //    sll x5 x11 x22      ====        sll t0, a1, s6
                                                  30'd    1884    : data = 32'h    C859CD93    ;    //    xori x27 x19 -891      ====        xori s11, s3, -891
                                                  30'd    1885    : data = 32'h    51AB7E13    ;    //    andi x28 x22 1306      ====        andi t3, s6, 1306
                                                  30'd    1886    : data = 32'h    80000937    ;    //    lui x18 524288      ====        li s2, 0x80000000 #start riscv_int_numeric_corner_stream_32
                                                  30'd    1887    : data = 32'h    00090913    ;    //    addi x18 x18 0      ====        li s2, 0x80000000 #start riscv_int_numeric_corner_stream_32
                                                  30'd    1888    : data = 32'h    0F77AC37    ;    //    lui x24 63354      ====        li s8, 0xf77987f
                                                  30'd    1889    : data = 32'h    87FC0C13    ;    //    addi x24 x24 -1921      ====        li s8, 0xf77987f
                                                  30'd    1890    : data = 32'h    00000993    ;    //    addi x19 x0 0      ====        li s3, 0x0
                                                  30'd    1891    : data = 32'h    80000EB7    ;    //    lui x29 524288      ====        li t4, 0x80000000
                                                  30'd    1892    : data = 32'h    000E8E93    ;    //    addi x29 x29 0      ====        li t4, 0x80000000
                                                  30'd    1893    : data = 32'h    7B8387B7    ;    //    lui x15 505912      ====        li a5, 0x7b83827a
                                                  30'd    1894    : data = 32'h    27A78793    ;    //    addi x15 x15 634      ====        li a5, 0x7b83827a
                                                  30'd    1895    : data = 32'h    00000F93    ;    //    addi x31 x0 0      ====        li t6, 0x0
                                                  30'd    1896    : data = 32'h    00000613    ;    //    addi x12 x0 0      ====        li a2, 0x0
                                                  30'd    1897    : data = 32'h    FFF00B13    ;    //    addi x22 x0 -1      ====        li s6, 0xffffffff
                                                  30'd    1898    : data = 32'h    00000893    ;    //    addi x17 x0 0      ====        li a7, 0x0
                                                  30'd    1899    : data = 32'h    A411CE37    ;    //    lui x28 672028      ====        li t3, 0xa411c375
                                                  30'd    1900    : data = 32'h    375E0E13    ;    //    addi x28 x28 885      ====        li t3, 0xa411c375
                                                  30'd    1901    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1902    : data = 32'h    418608B3    ;    //    sub x17 x12 x24      ====        sub a7, a2, s8
                                                  30'd    1903    : data = 32'h    41678B33    ;    //    sub x22 x15 x22      ====        sub s6, a5, s6
                                                  30'd    1904    : data = 32'h    41678633    ;    //    sub x12 x15 x22      ====        sub a2, a5, s6
                                                  30'd    1905    : data = 32'h    3BE5D797    ;    //    auipc x15 245341      ====        auipc a5, 245341
                                                  30'd    1906    : data = 32'h    41CE0B33    ;    //    sub x22 x28 x28      ====        sub s6, t3, t3
                                                  30'd    1907    : data = 32'h    4ED78793    ;    //    addi x15 x15 1261      ====        addi a5, a5, 1261
                                                  30'd    1908    : data = 32'h    01F90933    ;    //    add x18 x18 x31      ====        add s2, s2, t6
                                                  30'd    1909    : data = 32'h    995357B7    ;    //    lui x15 628021      ====        lui a5, 628021
                                                  30'd    1910    : data = 32'h    41CC0B33    ;    //    sub x22 x24 x28      ====        sub s6, s8, t3
                                                  30'd    1911    : data = 32'h    E2C287B7    ;    //    lui x15 928808      ====        lui a5, 928808
                                                  30'd    1912    : data = 32'h    CB378793    ;    //    addi x15 x15 -845      ====        addi a5, a5, -845
                                                  30'd    1913    : data = 32'h    ED641E97    ;    //    auipc x29 972353      ====        auipc t4, 972353
                                                  30'd    1914    : data = 32'h    EDE88613    ;    //    addi x12 x17 -290      ====        addi a2, a7, -290
                                                  30'd    1915    : data = 32'h    01DE0C33    ;    //    add x24 x28 x29      ====        add s8, t3, t4
                                                  30'd    1916    : data = 32'h    E32E8B13    ;    //    addi x22 x29 -462      ====        addi s6, t4, -462
                                                  30'd    1917    : data = 32'h    74B5D797    ;    //    auipc x15 478045      ====        auipc a5, 478045
                                                  30'd    1918    : data = 32'h    F32F8B13    ;    //    addi x22 x31 -206      ====        addi s6, t6, -206
                                                  30'd    1919    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1920    : data = 32'h    536E8893    ;    //    addi x17 x29 1334      ====        addi a7, t4, 1334
                                                  30'd    1921    : data = 32'h    01CB0FB3    ;    //    add x31 x22 x28      ====        add t6, s6, t3
                                                  30'd    1922    : data = 32'h    41688E33    ;    //    sub x28 x17 x22      ====        sub t3, a7, s6
                                                  30'd    1923    : data = 32'h    1DD95E17    ;    //    auipc x28 122261      ====        auipc t3, 122261
                                                  30'd    1924    : data = 32'h    B8133F97    ;    //    auipc x31 753971      ====        auipc t6, 753971
                                                  30'd    1925    : data = 32'h    B40B0913    ;    //    addi x18 x22 -1216      ====        addi s2, s6, -1216
                                                  30'd    1926    : data = 32'h    F9E60793    ;    //    addi x15 x12 -98      ====        addi a5, a2, -98
                                                  30'd    1927    : data = 32'h    41C787B3    ;    //    sub x15 x15 x28      ====        sub a5, a5, t3
                                                  30'd    1928    : data = 32'h    29AC0C13    ;    //    addi x24 x24 666      ====        addi s8, s8, 666
                                                  30'd    1929    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1930    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1931    : data = 32'h    0BD090EF    ;    //    jal x1 39100      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_32
                                                  30'd    1932    : data = 32'h    41DCDA33    ;    //    sra x20 x25 x29      ====        sra s4, s9, t4
                                                  30'd    1933    : data = 32'h    FB156593    ;    //    ori x11 x10 -79      ====        ori a1, a0, -79
                                                  30'd    1934    : data = 32'h    006B1813    ;    //    slli x16 x22 6      ====        slli a6, s6, 6
                                                  30'd    1935    : data = 32'h    B245A313    ;    //    slti x6 x11 -1244      ====        slti t1, a1, -1244
                                                  30'd    1936    : data = 32'h    001E0733    ;    //    add x14 x28 x1      ====        add a4, t3, ra
                                                  30'd    1937    : data = 32'h    41A48633    ;    //    sub x12 x9 x26      ====        sub a2, s1, s10
                                                  30'd    1938    : data = 32'h    016B58B3    ;    //    srl x17 x22 x22      ====        srl a7, s6, s6
                                                  30'd    1939    : data = 32'h    0010EB33    ;    //    or x22 x1 x1      ====        or s6, ra, ra
                                                  30'd    1940    : data = 32'h    95660037    ;    //    lui x0 611936      ====        lui zero, 611936
                                                  30'd    1941    : data = 32'h    00D90E33    ;    //    add x28 x18 x13      ====        add t3, s2, a3
                                                  30'd    1942    : data = 32'h    EAA2C413    ;    //    xori x8 x5 -342      ====        xori s0, t0, -342
                                                  30'd    1943    : data = 32'h    57F83813    ;    //    sltiu x16 x16 1407      ====        sltiu a6, a6, 1407
                                                  30'd    1944    : data = 32'h    7D70F893    ;    //    andi x17 x1 2007      ====        andi a7, ra, 2007
                                                  30'd    1945    : data = 32'h    005F9013    ;    //    slli x0 x31 5      ====        slli zero, t6, 5
                                                  30'd    1946    : data = 32'h    00325EB3    ;    //    srl x29 x4 x3      ====        srl t4, tp, gp
                                                  30'd    1947    : data = 32'h    0014CEB3    ;    //    xor x29 x9 x1      ====        xor t4, s1, ra
                                                  30'd    1948    : data = 32'h    41F10833    ;    //    sub x16 x2 x31      ====        sub a6, sp, t6
                                                  30'd    1949    : data = 32'h    80000C37    ;    //    lui x24 524288      ====        li s8, 0x80000000 #start riscv_int_numeric_corner_stream_11
                                                  30'd    1950    : data = 32'h    000C0C13    ;    //    addi x24 x24 0      ====        li s8, 0x80000000 #start riscv_int_numeric_corner_stream_11
                                                  30'd    1951    : data = 32'h    80000DB7    ;    //    lui x27 524288      ====        li s11, 0x80000000
                                                  30'd    1952    : data = 32'h    000D8D93    ;    //    addi x27 x27 0      ====        li s11, 0x80000000
                                                  30'd    1953    : data = 32'h    00000B93    ;    //    addi x23 x0 0      ====        li s7, 0x0
                                                  30'd    1954    : data = 32'h    368A99B7    ;    //    lui x19 223401      ====        li s3, 0x368a8f29
                                                  30'd    1955    : data = 32'h    F2998993    ;    //    addi x19 x19 -215      ====        li s3, 0x368a8f29
                                                  30'd    1956    : data = 32'h    FFF00493    ;    //    addi x9 x0 -1      ====        li s1, 0xffffffff
                                                  30'd    1957    : data = 32'h    50BE11B7    ;    //    lui x3 330721      ====        li gp, 0x50be0942
                                                  30'd    1958    : data = 32'h    94218193    ;    //    addi x3 x3 -1726      ====        li gp, 0x50be0942
                                                  30'd    1959    : data = 32'h    00000893    ;    //    addi x17 x0 0      ====        li a7, 0x0
                                                  30'd    1960    : data = 32'h    E6A5A937    ;    //    lui x18 944730      ====        li s2, 0xe6a5a304
                                                  30'd    1961    : data = 32'h    30490913    ;    //    addi x18 x18 772      ====        li s2, 0xe6a5a304
                                                  30'd    1962    : data = 32'h    00000A93    ;    //    addi x21 x0 0      ====        li s5, 0x0
                                                  30'd    1963    : data = 32'h    00000713    ;    //    addi x14 x0 0      ====        li a4, 0x0
                                                  30'd    1964    : data = 32'h    41298733    ;    //    sub x14 x19 x18      ====        sub a4, s3, s2
                                                  30'd    1965    : data = 32'h    403901B3    ;    //    sub x3 x18 x3      ====        sub gp, s2, gp
                                                  30'd    1966    : data = 32'h    CFC681B7    ;    //    lui x3 851048      ====        lui gp, 851048
                                                  30'd    1967    : data = 32'h    D6990C13    ;    //    addi x24 x18 -663      ====        addi s8, s2, -663
                                                  30'd    1968    : data = 32'h    6BA70A93    ;    //    addi x21 x14 1722      ====        addi s5, a4, 1722
                                                  30'd    1969    : data = 32'h    9D248D93    ;    //    addi x27 x9 -1582      ====        addi s11, s1, -1582
                                                  30'd    1970    : data = 32'h    018B8AB3    ;    //    add x21 x23 x24      ====        add s5, s7, s8
                                                  30'd    1971    : data = 32'h    BEA2B717    ;    //    auipc x14 780843      ====        auipc a4, 780843
                                                  30'd    1972    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1973    : data = 32'h    ACBB8C13    ;    //    addi x24 x23 -1333      ====        addi s8, s7, -1333
                                                  30'd    1974    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1975    : data = 32'h    017704B3    ;    //    add x9 x14 x23      ====        add s1, a4, s7
                                                  30'd    1976    : data = 32'h    017C08B3    ;    //    add x17 x24 x23      ====        add a7, s8, s7
                                                  30'd    1977    : data = 32'h    52C1E497    ;    //    auipc x9 338974      ====        auipc s1, 338974
                                                  30'd    1978    : data = 32'h    11D70913    ;    //    addi x18 x14 285      ====        addi s2, a4, 285
                                                  30'd    1979    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1980    : data = 32'h    939D8713    ;    //    addi x14 x27 -1735      ====        addi a4, s11, -1735
                                                  30'd    1981    : data = 32'h    D213AC17    ;    //    auipc x24 860474      ====        auipc s8, 860474
                                                  30'd    1982    : data = 32'h    40398733    ;    //    sub x14 x19 x3      ====        sub a4, s3, gp
                                                  30'd    1983    : data = 32'h    4FB5D717    ;    //    auipc x14 326493      ====        auipc a4, 326493
                                                  30'd    1984    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1985    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    1986    : data = 32'h    2EEB8713    ;    //    addi x14 x23 750      ====        addi a4, s7, 750
                                                  30'd    1987    : data = 32'h    41188933    ;    //    sub x18 x17 x17      ====        sub s2, a7, a7
                                                  30'd    1988    : data = 32'h    657E59B7    ;    //    lui x19 415717      ====        lui s3, 415717
                                                  30'd    1989    : data = 32'h    BCEDA8B7    ;    //    lui x17 773850      ====        lui a7, 773850
                                                  30'd    1990    : data = 32'h    949C7737    ;    //    lui x14 608711      ====        lui a4, 608711
                                                  30'd    1991    : data = 32'h    017A8C33    ;    //    add x24 x21 x23      ====        add s8, s5, s7
                                                  30'd    1992    : data = 32'h    01B98933    ;    //    add x18 x19 x27      ====        add s2, s3, s11
                                                  30'd    1993    : data = 32'h    7C4090EF    ;    //    jal x1 38852      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_11
                                                  30'd    1994    : data = 32'h    7A1BE113    ;    //    ori x2 x23 1953      ====        ori sp, s7, 1953
                                                  30'd    1995    : data = 32'h    C91DE413    ;    //    ori x8 x27 -879      ====        ori s0, s11, -879
                                                  30'd    1996    : data = 32'h    000717B3    ;    //    sll x15 x14 x0      ====        sll a5, a4, zero
                                                  30'd    1997    : data = 32'h    C3C5BE93    ;    //    sltiu x29 x11 -964      ====        sltiu t4, a1, -964
                                                  30'd    1998    : data = 32'h    0F8AB293    ;    //    sltiu x5 x21 248      ====        sltiu t0, s5, 248
                                                  30'd    1999    : data = 32'h    40DF0933    ;    //    sub x18 x30 x13      ====        sub s2, t5, a3
                                                  30'd    2000    : data = 32'h    E9280093    ;    //    addi x1 x16 -366      ====        addi ra, a6, -366
                                                  30'd    2001    : data = 32'h    019F34B3    ;    //    sltu x9 x30 x25      ====        sltu s1, t5, s9
                                                  30'd    2002    : data = 32'h    401A85B3    ;    //    sub x11 x21 x1      ====        sub a1, s5, ra
                                                  30'd    2003    : data = 32'h    3159F637    ;    //    lui x12 202143      ====        lui a2, 202143
                                                  30'd    2004    : data = 32'h    5524FA13    ;    //    andi x20 x9 1362      ====        andi s4, s1, 1362
                                                  30'd    2005    : data = 32'h    B9E5B017    ;    //    auipc x0 761435      ====        auipc zero, 761435
                                                  30'd    2006    : data = 32'h    0150DE93    ;    //    srli x29 x1 21      ====        srli t4, ra, 21
                                                  30'd    2007    : data = 32'h    2EE66593    ;    //    ori x11 x12 750      ====        ori a1, a2, 750
                                                  30'd    2008    : data = 32'h    33B50D93    ;    //    addi x27 x10 827      ====        addi s11, a0, 827
                                                  30'd    2009    : data = 32'h    00A11D13    ;    //    slli x26 x2 10      ====        slli s10, sp, 10
                                                  30'd    2010    : data = 32'h    001BBD33    ;    //    sltu x26 x23 x1      ====        sltu s10, s7, ra
                                                  30'd    2011    : data = 32'h    40108B33    ;    //    sub x22 x1 x1      ====        sub s6, ra, ra
                                                  30'd    2012    : data = 32'h    7B604837    ;    //    lui x16 505348      ====        lui a6, 505348
                                                  30'd    2013    : data = 32'h    14403793    ;    //    sltiu x15 x0 324      ====        sltiu a5, zero, 324
                                                  30'd    2014    : data = 32'h    8D22A597    ;    //    auipc x11 578090      ====        auipc a1, 578090
                                                  30'd    2015    : data = 32'h    40B85AB3    ;    //    sra x21 x16 x11      ====        sra s5, a6, a1
                                                  30'd    2016    : data = 32'h    AEEFA613    ;    //    slti x12 x31 -1298      ====        slti a2, t6, -1298
                                                  30'd    2017    : data = 32'h    01FA3333    ;    //    sltu x6 x20 x31      ====        sltu t1, s4, t6
                                                  30'd    2018    : data = 32'h    21A0F093    ;    //    andi x1 x1 538      ====        andi ra, ra, 538
                                                  30'd    2019    : data = 32'h    019C5D13    ;    //    srli x26 x24 25      ====        srli s10, s8, 25
                                                  30'd    2020    : data = 32'h    01249B33    ;    //    sll x22 x9 x18      ====        sll s6, s1, s2
                                                  30'd    2021    : data = 32'h    01351893    ;    //    slli x17 x10 19      ====        slli a7, a0, 19
                                                  30'd    2022    : data = 32'h    003DFB33    ;    //    and x22 x27 x3      ====        and s6, s11, gp
                                                  30'd    2023    : data = 32'h    40E7D0B3    ;    //    sra x1 x15 x14      ====        sra ra, a5, a4
                                                  30'd    2024    : data = 32'h    A41B3C13    ;    //    sltiu x24 x22 -1471      ====        sltiu s8, s6, -1471
                                                  30'd    2025    : data = 32'h    1EF76013    ;    //    ori x0 x14 495      ====        ori zero, a4, 495
                                                  30'd    2026    : data = 32'h    014CDA13    ;    //    srli x20 x25 20      ====        srli s4, s9, 20
                                                  30'd    2027    : data = 32'h    B2673C93    ;    //    sltiu x25 x14 -1242      ====        sltiu s9, a4, -1242
                                                  30'd    2028    : data = 32'h    00A3D493    ;    //    srli x9 x7 10      ====        srli s1, t2, 10
                                                  30'd    2029    : data = 32'h    4FC44A13    ;    //    xori x20 x8 1276      ====        xori s4, s0, 1276
                                                  30'd    2030    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2031    : data = 32'h    8A0C7293    ;    //    andi x5 x24 -1888      ====        andi t0, s8, -1888
                                                  30'd    2032    : data = 32'h    91C36C17    ;    //    auipc x24 597046      ====        auipc s8, 597046
                                                  30'd    2033    : data = 32'h    8B918413    ;    //    addi x8 x3 -1863      ====        addi s0, gp, -1863
                                                  30'd    2034    : data = 32'h    00B4C3B3    ;    //    xor x7 x9 x11      ====        xor t2, s1, a1
                                                  30'd    2035    : data = 32'h    00586333    ;    //    or x6 x16 x5      ====        or t1, a6, t0
                                                  30'd    2036    : data = 32'h    E529F913    ;    //    andi x18 x19 -430      ====        andi s2, s3, -430
                                                  30'd    2037    : data = 32'h    00FEDA93    ;    //    srli x21 x29 15      ====        srli s5, t4, 15
                                                  30'd    2038    : data = 32'h    4107D413    ;    //    srai x8 x15 16      ====        srai s0, a5, 16
                                                  30'd    2039    : data = 32'h    09B61DB7    ;    //    lui x27 39777      ====        lui s11, 39777
                                                  30'd    2040    : data = 32'h    017A3FB3    ;    //    sltu x31 x20 x23      ====        sltu t6, s4, s7
                                                  30'd    2041    : data = 32'h    C889F893    ;    //    andi x17 x19 -888      ====        andi a7, s3, -888
                                                  30'd    2042    : data = 32'h    00F29613    ;    //    slli x12 x5 15      ====        slli a2, t0, 15
                                                  30'd    2043    : data = 32'h    40640033    ;    //    sub x0 x8 x6      ====        sub zero, s0, t1
                                                  30'd    2044    : data = 32'h    AF2B4B93    ;    //    xori x23 x22 -1294      ====        xori s7, s6, -1294
                                                  30'd    2045    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2046    : data = 32'h    FBA78A13    ;    //    addi x20 x15 -70      ====        addi s4, a5, -70
                                                  30'd    2047    : data = 32'h    54A72B13    ;    //    slti x22 x14 1354      ====        slti s6, a4, 1354
                                                  30'd    2048    : data = 32'h    790F9437    ;    //    lui x8 495865      ====        lui s0, 495865
                                                  30'd    2049    : data = 32'h    2161A893    ;    //    slti x17 x3 534      ====        slti a7, gp, 534
                                                  30'd    2050    : data = 32'h    40000333    ;    //    sub x6 x0 x0      ====        sub t1, zero, zero
                                                  30'd    2051    : data = 32'h    804F7E17    ;    //    auipc x28 525559      ====        auipc t3, 525559
                                                  30'd    2052    : data = 32'h    50D7F013    ;    //    andi x0 x15 1293      ====        andi zero, a5, 1293
                                                  30'd    2053    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2054    : data = 32'h    B6398393    ;    //    addi x7 x19 -1181      ====        addi t2, s3, -1181
                                                  30'd    2055    : data = 32'h    0077A0B3    ;    //    slt x1 x15 x7      ====        slt ra, a5, t2
                                                  30'd    2056    : data = 32'h    5AE8F397    ;    //    auipc x7 372367      ====        auipc t2, 372367
                                                  30'd    2057    : data = 32'h    00465B13    ;    //    srli x22 x12 4      ====        srli s6, a2, 4
                                                  30'd    2058    : data = 32'h    95D435B7    ;    //    lui x11 613699      ====        lui a1, 613699
                                                  30'd    2059    : data = 32'h    0E16C693    ;    //    xori x13 x13 225      ====        xori a3, a3, 225
                                                  30'd    2060    : data = 32'h    00335893    ;    //    srli x17 x6 3      ====        srli a7, t1, 3
                                                  30'd    2061    : data = 32'h    40CEDB13    ;    //    srai x22 x29 12      ====        srai s6, t4, 12
                                                  30'd    2062    : data = 32'h    01FC5FB3    ;    //    srl x31 x24 x31      ====        srl t6, s8, t6
                                                  30'd    2063    : data = 32'h    0107EC33    ;    //    or x24 x15 x16      ====        or s8, a5, a6
                                                  30'd    2064    : data = 32'h    26D0F993    ;    //    andi x19 x1 621      ====        andi s3, ra, 621
                                                  30'd    2065    : data = 32'h    01835013    ;    //    srli x0 x6 24      ====        srli zero, t1, 24
                                                  30'd    2066    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2067    : data = 32'h    00271B13    ;    //    slli x22 x14 2      ====        slli s6, a4, 2
                                                  30'd    2068    : data = 32'h    003653B3    ;    //    srl x7 x12 x3      ====        srl t2, a2, gp
                                                  30'd    2069    : data = 32'h    862BCE93    ;    //    xori x29 x23 -1950      ====        xori t4, s7, -1950
                                                  30'd    2070    : data = 32'h    00633CB3    ;    //    sltu x25 x6 x6      ====        sltu s9, t1, t1
                                                  30'd    2071    : data = 32'h    CF7F5297    ;    //    auipc x5 849909      ====        auipc t0, 849909
                                                  30'd    2072    : data = 32'h    8EF02913    ;    //    slti x18 x0 -1809      ====        slti s2, zero, -1809
                                                  30'd    2073    : data = 32'h    0028EFB3    ;    //    or x31 x17 x2      ====        or t6, a7, sp
                                                  30'd    2074    : data = 32'h    35B34593    ;    //    xori x11 x6 859      ====        xori a1, t1, 859
                                                  30'd    2075    : data = 32'h    40B25813    ;    //    srai x16 x4 11      ====        srai a6, tp, 11
                                                  30'd    2076    : data = 32'h    5C69FA13    ;    //    andi x20 x19 1478      ====        andi s4, s3, 1478
                                                  30'd    2077    : data = 32'h    CEB13B37    ;    //    lui x22 846611      ====        lui s6, 846611
                                                  30'd    2078    : data = 32'h    BD5057B7    ;    //    lui x15 775429      ====        lui a5, 775429
                                                  30'd    2079    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2080    : data = 32'h    38118037    ;    //    lui x0 229656      ====        lui zero, 229656
                                                  30'd    2081    : data = 32'h    89A57413    ;    //    andi x8 x10 -1894      ====        andi s0, a0, -1894
                                                  30'd    2082    : data = 32'h    000BDA13    ;    //    srli x20 x23 0      ====        srli s4, s7, 0
                                                  30'd    2083    : data = 32'h    004837B3    ;    //    sltu x15 x16 x4      ====        sltu a5, a6, tp
                                                  30'd    2084    : data = 32'h    403E5A93    ;    //    srai x21 x28 3      ====        srai s5, t3, 3
                                                  30'd    2085    : data = 32'h    00A75D33    ;    //    srl x26 x14 x10      ====        srl s10, a4, a0
                                                  30'd    2086    : data = 32'h    40DD5CB3    ;    //    sra x25 x26 x13      ====        sra s9, s10, a3
                                                  30'd    2087    : data = 32'h    01C96B33    ;    //    or x22 x18 x28      ====        or s6, s2, t3
                                                  30'd    2088    : data = 32'h    5EA83C93    ;    //    sltiu x25 x16 1514      ====        sltiu s9, a6, 1514
                                                  30'd    2089    : data = 32'h    00825993    ;    //    srli x19 x4 8      ====        srli s3, tp, 8
                                                  30'd    2090    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2091    : data = 32'h    8448F893    ;    //    andi x17 x17 -1980      ====        andi a7, a7, -1980
                                                  30'd    2092    : data = 32'h    004CD6B3    ;    //    srl x13 x25 x4      ====        srl a3, s9, tp
                                                  30'd    2093    : data = 32'h    002FDB93    ;    //    srli x23 x31 2      ====        srli s7, t6, 2
                                                  30'd    2094    : data = 32'h    00BF7633    ;    //    and x12 x30 x11      ====        and a2, t5, a1
                                                  30'd    2095    : data = 32'h    403DD0B3    ;    //    sra x1 x27 x3      ====        sra ra, s11, gp
                                                  30'd    2096    : data = 32'h    408BD2B3    ;    //    sra x5 x23 x8      ====        sra t0, s7, s0
                                                  30'd    2097    : data = 32'h    C3D4C793    ;    //    xori x15 x9 -963      ====        xori a5, s1, -963
                                                  30'd    2098    : data = 32'h    01287433    ;    //    and x8 x16 x18      ====        and s0, a6, s2
                                                  30'd    2099    : data = 32'h    01934033    ;    //    xor x0 x6 x25      ====        xor zero, t1, s9
                                                  30'd    2100    : data = 32'h    66EC6CB7    ;    //    lui x25 421574      ====        lui s9, 421574
                                                  30'd    2101    : data = 32'h    41192A93    ;    //    slti x21 x18 1041      ====        slti s5, s2, 1041
                                                  30'd    2102    : data = 32'h    F0AB8613    ;    //    addi x12 x23 -246      ====        addi a2, s7, -246
                                                  30'd    2103    : data = 32'h    01F186B3    ;    //    add x13 x3 x31      ====        add a3, gp, t6
                                                  30'd    2104    : data = 32'h    0932F893    ;    //    andi x17 x5 147      ====        andi a7, t0, 147
                                                  30'd    2105    : data = 32'h    31F0C413    ;    //    xori x8 x1 799      ====        xori s0, ra, 799
                                                  30'd    2106    : data = 32'h    009B6CB3    ;    //    or x25 x22 x9      ====        or s9, s6, s1
                                                  30'd    2107    : data = 32'h    C5397793    ;    //    andi x15 x18 -941      ====        andi a5, s2, -941
                                                  30'd    2108    : data = 32'h    0036D613    ;    //    srli x12 x13 3      ====        srli a2, a3, 3
                                                  30'd    2109    : data = 32'h    01ECAB33    ;    //    slt x22 x25 x30      ====        slt s6, s9, t5
                                                  30'd    2110    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2111    : data = 32'h    406759B3    ;    //    sra x19 x14 x6      ====        sra s3, a4, t1
                                                  30'd    2112    : data = 32'h    013D9C13    ;    //    slli x24 x27 19      ====        slli s8, s11, 19
                                                  30'd    2113    : data = 32'h    40930933    ;    //    sub x18 x6 x9      ====        sub s2, t1, s1
                                                  30'd    2114    : data = 32'h    C574CE13    ;    //    xori x28 x9 -937      ====        xori t3, s1, -937
                                                  30'd    2115    : data = 32'h    010F1B93    ;    //    slli x23 x30 16      ====        slli s7, t5, 16
                                                  30'd    2116    : data = 32'h    41085EB3    ;    //    sra x29 x16 x16      ====        sra t4, a6, a6
                                                  30'd    2117    : data = 32'h    2A0A7B13    ;    //    andi x22 x20 672      ====        andi s6, s4, 672
                                                  30'd    2118    : data = 32'h    4157D013    ;    //    srai x0 x15 21      ====        srai zero, a5, 21
                                                  30'd    2119    : data = 32'h    0162AEB3    ;    //    slt x29 x5 x22      ====        slt t4, t0, s6
                                                  30'd    2120    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2121    : data = 32'h    00D208B3    ;    //    add x17 x4 x13      ====        add a7, tp, a3
                                                  30'd    2122    : data = 32'h    00568D33    ;    //    add x26 x13 x5      ====        add s10, a3, t0
                                                  30'd    2123    : data = 32'h    411ED2B3    ;    //    sra x5 x29 x17      ====        sra t0, t4, a7
                                                  30'd    2124    : data = 32'h    0033DD93    ;    //    srli x27 x7 3      ====        srli s11, t2, 3
                                                  30'd    2125    : data = 32'h    01894D33    ;    //    xor x26 x18 x24      ====        xor s10, s2, s8
                                                  30'd    2126    : data = 32'h    2F94AE93    ;    //    slti x29 x9 761      ====        slti t4, s1, 761
                                                  30'd    2127    : data = 32'h    01969713    ;    //    slli x14 x13 25      ====        slli a4, a3, 25
                                                  30'd    2128    : data = 32'h    A761BC13    ;    //    sltiu x24 x3 -1418      ====        sltiu s8, gp, -1418
                                                  30'd    2129    : data = 32'h    FBB0FE13    ;    //    andi x28 x1 -69      ====        andi t3, ra, -69
                                                  30'd    2130    : data = 32'h    01378DB3    ;    //    add x27 x15 x19      ====        add s11, a5, s3
                                                  30'd    2131    : data = 32'h    00B79C13    ;    //    slli x24 x15 11      ====        slli s8, a5, 11
                                                  30'd    2132    : data = 32'h    00EF9A93    ;    //    slli x21 x31 14      ====        slli s5, t6, 14
                                                  30'd    2133    : data = 32'h    123F5CB7    ;    //    lui x25 74741      ====        lui s9, 74741
                                                  30'd    2134    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2135    : data = 32'h    0125DA13    ;    //    srli x20 x11 18      ====        srli s4, a1, 18
                                                  30'd    2136    : data = 32'h    005D0733    ;    //    add x14 x26 x5      ====        add a4, s10, t0
                                                  30'd    2137    : data = 32'h    0123BFB3    ;    //    sltu x31 x7 x18      ====        sltu t6, t2, s2
                                                  30'd    2138    : data = 32'h    402ED5B3    ;    //    sra x11 x29 x2      ====        sra a1, t4, sp
                                                  30'd    2139    : data = 32'h    1D534293    ;    //    xori x5 x6 469      ====        xori t0, t1, 469
                                                  30'd    2140    : data = 32'h    002E9393    ;    //    slli x7 x29 2      ====        slli t2, t4, 2
                                                  30'd    2141    : data = 32'h    D011B893    ;    //    sltiu x17 x3 -767      ====        sltiu a7, gp, -767
                                                  30'd    2142    : data = 32'h    89B4CC17    ;    //    auipc x24 564044      ====        auipc s8, 564044
                                                  30'd    2143    : data = 32'h    0E1ECC97    ;    //    auipc x25 57836      ====        auipc s9, 57836
                                                  30'd    2144    : data = 32'h    3CD04417    ;    //    auipc x8 249092      ====        auipc s0, 249092
                                                  30'd    2145    : data = 32'h    2DB459B7    ;    //    lui x19 187205      ====        lui s3, 187205
                                                  30'd    2146    : data = 32'h    40FC5E13    ;    //    srai x28 x24 15      ====        srai t3, s8, 15
                                                  30'd    2147    : data = 32'h    C97DAFB7    ;    //    lui x31 825306      ====        lui t6, 825306
                                                  30'd    2148    : data = 32'h    01DF28B3    ;    //    slt x17 x30 x29      ====        slt a7, t5, t4
                                                  30'd    2149    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2150    : data = 32'h    018626B3    ;    //    slt x13 x12 x24      ====        slt a3, a2, s8
                                                  30'd    2151    : data = 32'h    D7BBB013    ;    //    sltiu x0 x23 -645      ====        sltiu zero, s7, -645
                                                  30'd    2152    : data = 32'h    2EEB3593    ;    //    sltiu x11 x22 750      ====        sltiu a1, s6, 750
                                                  30'd    2153    : data = 32'h    5DCA0F93    ;    //    addi x31 x20 1500      ====        addi t6, s4, 1500
                                                  30'd    2154    : data = 32'h    0032D3B3    ;    //    srl x7 x5 x3      ====        srl t2, t0, gp
                                                  30'd    2155    : data = 32'h    23A7E193    ;    //    ori x3 x15 570      ====        ori gp, a5, 570
                                                  30'd    2156    : data = 32'h    01CF2E33    ;    //    slt x28 x30 x28      ====        slt t3, t5, t3
                                                  30'd    2157    : data = 32'h    413DDD33    ;    //    sra x26 x27 x19      ====        sra s10, s11, s3
                                                  30'd    2158    : data = 32'h    0016C733    ;    //    xor x14 x13 x1      ====        xor a4, a3, ra
                                                  30'd    2159    : data = 32'h    116F0113    ;    //    addi x2 x30 278      ====        addi sp, t5, 278
                                                  30'd    2160    : data = 32'h    01F2D733    ;    //    srl x14 x5 x31      ====        srl a4, t0, t6
                                                  30'd    2161    : data = 32'h    41755B13    ;    //    srai x22 x10 23      ====        srai s6, a0, 23
                                                  30'd    2162    : data = 32'h    40A5D6B3    ;    //    sra x13 x11 x10      ====        sra a3, a1, a0
                                                  30'd    2163    : data = 32'h    98A6B493    ;    //    sltiu x9 x13 -1654      ====        sltiu s1, a3, -1654
                                                  30'd    2164    : data = 32'h    5193E813    ;    //    ori x16 x7 1305      ====        ori a6, t2, 1305
                                                  30'd    2165    : data = 32'h    FC8E6C93    ;    //    ori x25 x28 -56      ====        ori s9, t3, -56
                                                  30'd    2166    : data = 32'h    0142C933    ;    //    xor x18 x5 x20      ====        xor s2, t0, s4
                                                  30'd    2167    : data = 32'h    98552B13    ;    //    slti x22 x10 -1659      ====        slti s6, a0, -1659
                                                  30'd    2168    : data = 32'h    FF84CF93    ;    //    xori x31 x9 -8      ====        xori t6, s1, -8
                                                  30'd    2169    : data = 32'h    01AF5BB3    ;    //    srl x23 x30 x26      ====        srl s7, t5, s10
                                                  30'd    2170    : data = 32'h    0C6EECB7    ;    //    lui x25 50926      ====        lui s9, 50926
                                                  30'd    2171    : data = 32'h    415B8BB3    ;    //    sub x23 x23 x21      ====        sub s7, s7, s5
                                                  30'd    2172    : data = 32'h    997923B7    ;    //    lui x7 628626      ====        lui t2, 628626
                                                  30'd    2173    : data = 32'h    40E38633    ;    //    sub x12 x7 x14      ====        sub a2, t2, a4
                                                  30'd    2174    : data = 32'h    A8216A93    ;    //    ori x21 x2 -1406      ====        ori s5, sp, -1406
                                                  30'd    2175    : data = 32'h    A0CA6093    ;    //    ori x1 x20 -1524      ====        ori ra, s4, -1524
                                                  30'd    2176    : data = 32'h    41E35713    ;    //    srai x14 x6 30      ====        srai a4, t1, 30
                                                  30'd    2177    : data = 32'h    01859413    ;    //    slli x8 x11 24      ====        slli s0, a1, 24
                                                  30'd    2178    : data = 32'h    4404A293    ;    //    slti x5 x9 1088      ====        slti t0, s1, 1088
                                                  30'd    2179    : data = 32'h    BE320317    ;    //    auipc x6 779040      ====        auipc t1, 779040
                                                  30'd    2180    : data = 32'h    40A9D133    ;    //    sra x2 x19 x10      ====        sra sp, s3, a0
                                                  30'd    2181    : data = 32'h    0109B433    ;    //    sltu x8 x19 x16      ====        sltu s0, s3, a6
                                                  30'd    2182    : data = 32'h    0176A633    ;    //    slt x12 x13 x23      ====        slt a2, a3, s7
                                                  30'd    2183    : data = 32'h    00F066B3    ;    //    or x13 x0 x15      ====        or a3, zero, a5
                                                  30'd    2184    : data = 32'h    051E7693    ;    //    andi x13 x28 81      ====        andi a3, t3, 81
                                                  30'd    2185    : data = 32'h    89F4AC13    ;    //    slti x24 x9 -1889      ====        slti s8, s1, -1889
                                                  30'd    2186    : data = 32'h    40910333    ;    //    sub x6 x2 x9      ====        sub t1, sp, s1
                                                  30'd    2187    : data = 32'h    41B45B33    ;    //    sra x22 x8 x27      ====        sra s6, s0, s11
                                                  30'd    2188    : data = 32'h    CC9B4A13    ;    //    xori x20 x22 -823      ====        xori s4, s6, -823
                                                  30'd    2189    : data = 32'h    A0646893    ;    //    ori x17 x8 -1530      ====        ori a7, s0, -1530
                                                  30'd    2190    : data = 32'h    01E281B3    ;    //    add x3 x5 x30      ====        add gp, t0, t5
                                                  30'd    2191    : data = 32'h    406ADC13    ;    //    srai x24 x21 6      ====        srai s8, s5, 6
                                                  30'd    2192    : data = 32'h    002242B3    ;    //    xor x5 x4 x2      ====        xor t0, tp, sp
                                                  30'd    2193    : data = 32'h    00924E33    ;    //    xor x28 x4 x9      ====        xor t3, tp, s1
                                                  30'd    2194    : data = 32'h    01B7D6B3    ;    //    srl x13 x15 x27      ====        srl a3, a5, s11
                                                  30'd    2195    : data = 32'h    01B17A33    ;    //    and x20 x2 x27      ====        and s4, sp, s11
                                                  30'd    2196    : data = 32'h    A2787C37    ;    //    lui x24 665479      ====        lui s8, 665479
                                                  30'd    2197    : data = 32'h    00C040B3    ;    //    xor x1 x0 x12      ====        xor ra, zero, a2
                                                  30'd    2198    : data = 32'h    007107B3    ;    //    add x15 x2 x7      ====        add a5, sp, t2
                                                  30'd    2199    : data = 32'h    0135D293    ;    //    srli x5 x11 19      ====        srli t0, a1, 19
                                                  30'd    2200    : data = 32'h    0010A2B3    ;    //    slt x5 x1 x1      ====        slt t0, ra, ra
                                                  30'd    2201    : data = 32'h    0034D5B3    ;    //    srl x11 x9 x3      ====        srl a1, s1, gp
                                                  30'd    2202    : data = 32'h    41DF89B3    ;    //    sub x19 x31 x29      ====        sub s3, t6, t4
                                                  30'd    2203    : data = 32'h    0026D2B3    ;    //    srl x5 x13 x2      ====        srl t0, a3, sp
                                                  30'd    2204    : data = 32'h    A62801B7    ;    //    lui x3 680576      ====        lui gp, 680576
                                                  30'd    2205    : data = 32'h    019DE133    ;    //    or x2 x27 x25      ====        or sp, s11, s9
                                                  30'd    2206    : data = 32'h    01495C13    ;    //    srli x24 x18 20      ====        srli s8, s2, 20
                                                  30'd    2207    : data = 32'h    D0EE50B7    ;    //    lui x1 855781      ====        lui ra, 855781
                                                  30'd    2208    : data = 32'h    012E1B13    ;    //    slli x22 x28 18      ====        slli s6, t3, 18
                                                  30'd    2209    : data = 32'h    95B4BA93    ;    //    sltiu x21 x9 -1701      ====        sltiu s5, s1, -1701
                                                  30'd    2210    : data = 32'h    013FF933    ;    //    and x18 x31 x19      ====        and s2, t6, s3
                                                  30'd    2211    : data = 32'h    015A57B3    ;    //    srl x15 x20 x21      ====        srl a5, s4, s5
                                                  30'd    2212    : data = 32'h    8DF236B7    ;    //    lui x13 581411      ====        lui a3, 581411
                                                  30'd    2213    : data = 32'h    41C4DB33    ;    //    sra x22 x9 x28      ====        sra s6, s1, t3
                                                  30'd    2214    : data = 32'h    012085B3    ;    //    add x11 x1 x18      ====        add a1, ra, s2
                                                  30'd    2215    : data = 32'h    4F2A7F93    ;    //    andi x31 x20 1266      ====        andi t6, s4, 1266
                                                  30'd    2216    : data = 32'h    00F55B33    ;    //    srl x22 x10 x15      ====        srl s6, a0, a5
                                                  30'd    2217    : data = 32'h    004FD8B3    ;    //    srl x17 x31 x4      ====        srl a7, t6, tp
                                                  30'd    2218    : data = 32'h    407185B3    ;    //    sub x11 x3 x7      ====        sub a1, gp, t2
                                                  30'd    2219    : data = 32'h    01786E33    ;    //    or x28 x16 x23      ====        or t3, a6, s7
                                                  30'd    2220    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2221    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2222    : data = 32'h    00C375B3    ;    //    and x11 x6 x12      ====        and a1, t1, a2
                                                  30'd    2223    : data = 32'h    D62BE117    ;    //    auipc x2 877246      ====        auipc sp, 877246
                                                  30'd    2224    : data = 32'h    00A76D33    ;    //    or x26 x14 x10      ====        or s10, a4, a0
                                                  30'd    2225    : data = 32'h    254F6DB7    ;    //    lui x27 152822      ====        lui s11, 152822
                                                  30'd    2226    : data = 32'h    00E81A13    ;    //    slli x20 x16 14      ====        slli s4, a6, 14
                                                  30'd    2227    : data = 32'h    410A5013    ;    //    srai x0 x20 16      ====        srai zero, s4, 16
                                                  30'd    2228    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2229    : data = 32'h    A1022E93    ;    //    slti x29 x4 -1520      ====        slti t4, tp, -1520
                                                  30'd    2230    : data = 32'h    40B60D33    ;    //    sub x26 x12 x11      ====        sub s10, a2, a1
                                                  30'd    2231    : data = 32'h    006F9933    ;    //    sll x18 x31 x6      ====        sll s2, t6, t1
                                                  30'd    2232    : data = 32'h    4366E713    ;    //    ori x14 x13 1078      ====        ori a4, a3, 1078
                                                  30'd    2233    : data = 32'h    96E20693    ;    //    addi x13 x4 -1682      ====        addi a3, tp, -1682
                                                  30'd    2234    : data = 32'h    01553AB3    ;    //    sltu x21 x10 x21      ====        sltu s5, a0, s5
                                                  30'd    2235    : data = 32'h    1E09F493    ;    //    andi x9 x19 480      ====        andi s1, s3, 480
                                                  30'd    2236    : data = 32'h    016F1E93    ;    //    slli x29 x30 22      ====        slli t4, t5, 22
                                                  30'd    2237    : data = 32'h    2860F613    ;    //    andi x12 x1 646      ====        andi a2, ra, 646
                                                  30'd    2238    : data = 32'h    00085A13    ;    //    srli x20 x16 0      ====        srli s4, a6, 0
                                                  30'd    2239    : data = 32'h    00B7BFB3    ;    //    sltu x31 x15 x11      ====        sltu t6, a5, a1
                                                  30'd    2240    : data = 32'h    4E1BCC13    ;    //    xori x24 x23 1249      ====        xori s8, s7, 1249
                                                  30'd    2241    : data = 32'h    01DC20B3    ;    //    slt x1 x24 x29      ====        slt ra, s8, t4
                                                  30'd    2242    : data = 32'h    016BDD13    ;    //    srli x26 x23 22      ====        srli s10, s7, 22
                                                  30'd    2243    : data = 32'h    0145F1B3    ;    //    and x3 x11 x20      ====        and gp, a1, s4
                                                  30'd    2244    : data = 32'h    41C85FB3    ;    //    sra x31 x16 x28      ====        sra t6, a6, t3
                                                  30'd    2245    : data = 32'h    4133DB93    ;    //    srai x23 x7 19      ====        srai s7, t2, 19
                                                  30'd    2246    : data = 32'h    00791933    ;    //    sll x18 x18 x7      ====        sll s2, s2, t2
                                                  30'd    2247    : data = 32'h    00594D33    ;    //    xor x26 x18 x5      ====        xor s10, s2, t0
                                                  30'd    2248    : data = 32'h    0022AFB3    ;    //    slt x31 x5 x2      ====        slt t6, t0, sp
                                                  30'd    2249    : data = 32'h    01C18E33    ;    //    add x28 x3 x28      ====        add t3, gp, t3
                                                  30'd    2250    : data = 32'h    00FFE733    ;    //    or x14 x31 x15      ====        or a4, t6, a5
                                                  30'd    2251    : data = 32'h    01D6AE33    ;    //    slt x28 x13 x29      ====        slt t3, a3, t4
                                                  30'd    2252    : data = 32'h    00566033    ;    //    or x0 x12 x5      ====        or zero, a2, t0
                                                  30'd    2253    : data = 32'h    8ED14713    ;    //    xori x14 x2 -1811      ====        xori a4, sp, -1811
                                                  30'd    2254    : data = 32'h    8B246397    ;    //    auipc x7 569926      ====        auipc t2, 569926
                                                  30'd    2255    : data = 32'h    00E6CD33    ;    //    xor x26 x13 x14      ====        xor s10, a3, a4
                                                  30'd    2256    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2257    : data = 32'h    00F879B3    ;    //    and x19 x16 x15      ====        and s3, a6, a5
                                                  30'd    2258    : data = 32'h    A381C013    ;    //    xori x0 x3 -1480      ====        xori zero, gp, -1480
                                                  30'd    2259    : data = 32'h    30E5E013    ;    //    ori x0 x11 782      ====        ori zero, a1, 782
                                                  30'd    2260    : data = 32'h    339C3193    ;    //    sltiu x3 x24 825      ====        sltiu gp, s8, 825
                                                  30'd    2261    : data = 32'h    A233E913    ;    //    ori x18 x7 -1501      ====        ori s2, t2, -1501
                                                  30'd    2262    : data = 32'h    008A2BB3    ;    //    slt x23 x20 x8      ====        slt s7, s4, s0
                                                  30'd    2263    : data = 32'h    0B3CCD37    ;    //    lui x26 46028      ====        lui s10, 46028
                                                  30'd    2264    : data = 32'h    01501613    ;    //    slli x12 x0 21      ====        slli a2, zero, 21
                                                  30'd    2265    : data = 32'h    00FECBB3    ;    //    xor x23 x29 x15      ====        xor s7, t4, a5
                                                  30'd    2266    : data = 32'h    004F8733    ;    //    add x14 x31 x4      ====        add a4, t6, tp
                                                  30'd    2267    : data = 32'h    01EC1793    ;    //    slli x15 x24 30      ====        slli a5, s8, 30
                                                  30'd    2268    : data = 32'h    004C5A93    ;    //    srli x21 x24 4      ====        srli s5, s8, 4
                                                  30'd    2269    : data = 32'h    3FF92A13    ;    //    slti x20 x18 1023      ====        slti s4, s2, 1023
                                                  30'd    2270    : data = 32'h    01B1F2B3    ;    //    and x5 x3 x27      ====        and t0, gp, s11
                                                  30'd    2271    : data = 32'h    016DE5B3    ;    //    or x11 x27 x22      ====        or a1, s11, s6
                                                  30'd    2272    : data = 32'h    011CDC33    ;    //    srl x24 x25 x17      ====        srl s8, s9, a7
                                                  30'd    2273    : data = 32'h    43509497    ;    //    auipc x9 275721      ====        auipc s1, 275721
                                                  30'd    2274    : data = 32'h    00354633    ;    //    xor x12 x10 x3      ====        xor a2, a0, gp
                                                  30'd    2275    : data = 32'h    2190E593    ;    //    ori x11 x1 537      ====        ori a1, ra, 537
                                                  30'd    2276    : data = 32'h    003C8B33    ;    //    add x22 x25 x3      ====        add s6, s9, gp
                                                  30'd    2277    : data = 32'h    01D28433    ;    //    add x8 x5 x29      ====        add s0, t0, t4
                                                  30'd    2278    : data = 32'h    002D3033    ;    //    sltu x0 x26 x2      ====        sltu zero, s10, sp
                                                  30'd    2279    : data = 32'h    01AFF3B3    ;    //    and x7 x31 x26      ====        and t2, t6, s10
                                                  30'd    2280    : data = 32'h    88E0BB13    ;    //    sltiu x22 x1 -1906      ====        sltiu s6, ra, -1906
                                                  30'd    2281    : data = 32'h    003D32B3    ;    //    sltu x5 x26 x3      ====        sltu t0, s10, gp
                                                  30'd    2282    : data = 32'h    40740633    ;    //    sub x12 x8 x7      ====        sub a2, s0, t2
                                                  30'd    2283    : data = 32'h    00A67133    ;    //    and x2 x12 x10      ====        and sp, a2, a0
                                                  30'd    2284    : data = 32'h    00CF1293    ;    //    slli x5 x30 12      ====        slli t0, t5, 12
                                                  30'd    2285    : data = 32'h    01E69813    ;    //    slli x16 x13 30      ====        slli a6, a3, 30
                                                  30'd    2286    : data = 32'h    AC6A9917    ;    //    auipc x18 706217      ====        auipc s2, 706217
                                                  30'd    2287    : data = 32'h    0049D0B3    ;    //    srl x1 x19 x4      ====        srl ra, s3, tp
                                                  30'd    2288    : data = 32'h    01E71133    ;    //    sll x2 x14 x30      ====        sll sp, a4, t5
                                                  30'd    2289    : data = 32'h    01EB9AB3    ;    //    sll x21 x23 x30      ====        sll s5, s7, t5
                                                  30'd    2290    : data = 32'h    C2377913    ;    //    andi x18 x14 -989      ====        andi s2, a4, -989
                                                  30'd    2291    : data = 32'h    003AA0B3    ;    //    slt x1 x21 x3      ====        slt ra, s5, gp
                                                  30'd    2292    : data = 32'h    14F43A93    ;    //    sltiu x21 x8 335      ====        sltiu s5, s0, 335
                                                  30'd    2293    : data = 32'h    01CAF6B3    ;    //    and x13 x21 x28      ====        and a3, s5, t3
                                                  30'd    2294    : data = 32'h    01CC1593    ;    //    slli x11 x24 28      ====        slli a1, s8, 28
                                                  30'd    2295    : data = 32'h    00786133    ;    //    or x2 x16 x7      ====        or sp, a6, t2
                                                  30'd    2296    : data = 32'h    00259DB3    ;    //    sll x27 x11 x2      ====        sll s11, a1, sp
                                                  30'd    2297    : data = 32'h    00E0C3B3    ;    //    xor x7 x1 x14      ====        xor t2, ra, a4
                                                  30'd    2298    : data = 32'h    0176BD33    ;    //    sltu x26 x13 x23      ====        sltu s10, a3, s7
                                                  30'd    2299    : data = 32'h    08A7EA93    ;    //    ori x21 x15 138      ====        ori s5, a5, 138
                                                  30'd    2300    : data = 32'h    13B9F293    ;    //    andi x5 x19 315      ====        andi t0, s3, 315
                                                  30'd    2301    : data = 32'h    8FCAAB93    ;    //    slti x23 x21 -1796      ====        slti s7, s5, -1796
                                                  30'd    2302    : data = 32'h    40CF5313    ;    //    srai x6 x30 12      ====        srai t1, t5, 12
                                                  30'd    2303    : data = 32'h    003ED093    ;    //    srli x1 x29 3      ====        srli ra, t4, 3
                                                  30'd    2304    : data = 32'h    403ED813    ;    //    srai x16 x29 3      ====        srai a6, t4, 3
                                                  30'd    2305    : data = 32'h    9A5A0C93    ;    //    addi x25 x20 -1627      ====        addi s9, s4, -1627
                                                  30'd    2306    : data = 32'h    00D4E5B3    ;    //    or x11 x9 x13      ====        or a1, s1, a3
                                                  30'd    2307    : data = 32'h    0031F633    ;    //    and x12 x3 x3      ====        and a2, gp, gp
                                                  30'd    2308    : data = 32'h    B2765A97    ;    //    auipc x21 730981      ====        auipc s5, 730981
                                                  30'd    2309    : data = 32'h    40CF84B3    ;    //    sub x9 x31 x12      ====        sub s1, t6, a2
                                                  30'd    2310    : data = 32'h    00111193    ;    //    slli x3 x2 1      ====        slli gp, sp, 1
                                                  30'd    2311    : data = 32'h    91B72413    ;    //    slti x8 x14 -1765      ====        slti s0, a4, -1765
                                                  30'd    2312    : data = 32'h    CAE0B437    ;    //    lui x8 830987      ====        lui s0, 830987
                                                  30'd    2313    : data = 32'h    010E2933    ;    //    slt x18 x28 x16      ====        slt s2, t3, a6
                                                  30'd    2314    : data = 32'h    36428937    ;    //    lui x18 222248      ====        lui s2, 222248
                                                  30'd    2315    : data = 32'h    00B88133    ;    //    add x2 x17 x11      ====        add sp, a7, a1
                                                  30'd    2316    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2317    : data = 32'h    00B51393    ;    //    slli x7 x10 11      ====        slli t2, a0, 11
                                                  30'd    2318    : data = 32'h    000749B3    ;    //    xor x19 x14 x0      ====        xor s3, a4, zero
                                                  30'd    2319    : data = 32'h    40F9DBB3    ;    //    sra x23 x19 x15      ====        sra s7, s3, a5
                                                  30'd    2320    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2321    : data = 32'h    B6D58713    ;    //    addi x14 x11 -1171      ====        addi a4, a1, -1171
                                                  30'd    2322    : data = 32'h    01A6D293    ;    //    srli x5 x13 26      ====        srli t0, a3, 26
                                                  30'd    2323    : data = 32'h    A51CD697    ;    //    auipc x13 676301      ====        auipc a3, 676301
                                                  30'd    2324    : data = 32'h    E4BC0713    ;    //    addi x14 x24 -437      ====        addi a4, s8, -437
                                                  30'd    2325    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2326    : data = 32'h    01C05EB3    ;    //    srl x29 x0 x28      ====        srl t4, zero, t3
                                                  30'd    2327    : data = 32'h    C6864193    ;    //    xori x3 x12 -920      ====        xori gp, a2, -920
                                                  30'd    2328    : data = 32'h    40A7DD93    ;    //    srai x27 x15 10      ====        srai s11, a5, 10
                                                  30'd    2329    : data = 32'h    41FB8633    ;    //    sub x12 x23 x31      ====        sub a2, s7, t6
                                                  30'd    2330    : data = 32'h    40F15A13    ;    //    srai x20 x2 15      ====        srai s4, sp, 15
                                                  30'd    2331    : data = 32'h    E2793C13    ;    //    sltiu x24 x18 -473      ====        sltiu s8, s2, -473
                                                  30'd    2332    : data = 32'h    DEAF7B13    ;    //    andi x22 x30 -534      ====        andi s6, t5, -534
                                                  30'd    2333    : data = 32'h    60352613    ;    //    slti x12 x10 1539      ====        slti a2, a0, 1539
                                                  30'd    2334    : data = 32'h    8A3EF813    ;    //    andi x16 x29 -1885      ====        andi a6, t4, -1885
                                                  30'd    2335    : data = 32'h    01B97BB3    ;    //    and x23 x18 x27      ====        and s7, s2, s11
                                                  30'd    2336    : data = 32'h    410C8933    ;    //    sub x18 x25 x16      ====        sub s2, s9, a6
                                                  30'd    2337    : data = 32'h    41475033    ;    //    sra x0 x14 x20      ====        sra zero, a4, s4
                                                  30'd    2338    : data = 32'h    F1A04BB7    ;    //    lui x23 989700      ====        lui s7, 989700
                                                  30'd    2339    : data = 32'h    4145D993    ;    //    srai x19 x11 20      ====        srai s3, a1, 20
                                                  30'd    2340    : data = 32'h    408587B3    ;    //    sub x15 x11 x8      ====        sub a5, a1, s0
                                                  30'd    2341    : data = 32'h    016DFAB3    ;    //    and x21 x27 x22      ====        and s5, s11, s6
                                                  30'd    2342    : data = 32'h    E69CE713    ;    //    ori x14 x25 -407      ====        ori a4, s9, -407
                                                  30'd    2343    : data = 32'h    649A7593    ;    //    andi x11 x20 1609      ====        andi a1, s4, 1609
                                                  30'd    2344    : data = 32'h    0175F133    ;    //    and x2 x11 x23      ====        and sp, a1, s7
                                                  30'd    2345    : data = 32'h    9B4BB613    ;    //    sltiu x12 x23 -1612      ====        sltiu a2, s7, -1612
                                                  30'd    2346    : data = 32'h    00DD5D33    ;    //    srl x26 x26 x13      ====        srl s10, s10, a3
                                                  30'd    2347    : data = 32'h    0074D033    ;    //    srl x0 x9 x7      ====        srl zero, s1, t2
                                                  30'd    2348    : data = 32'h    004A55B3    ;    //    srl x11 x20 x4      ====        srl a1, s4, tp
                                                  30'd    2349    : data = 32'h    2723CB93    ;    //    xori x23 x7 626      ====        xori s7, t2, 626
                                                  30'd    2350    : data = 32'h    CA2598B7    ;    //    lui x17 827993      ====        lui a7, 827993
                                                  30'd    2351    : data = 32'h    015C6733    ;    //    or x14 x24 x21      ====        or a4, s8, s5
                                                  30'd    2352    : data = 32'h    01930B33    ;    //    add x22 x6 x25      ====        add s6, t1, s9
                                                  30'd    2353    : data = 32'h    41188C33    ;    //    sub x24 x17 x17      ====        sub s8, a7, a7
                                                  30'd    2354    : data = 32'h    831DCD13    ;    //    xori x26 x27 -1999      ====        xori s10, s11, -1999
                                                  30'd    2355    : data = 32'h    0004E433    ;    //    or x8 x9 x0      ====        or s0, s1, zero
                                                  30'd    2356    : data = 32'h    001BDB33    ;    //    srl x22 x23 x1      ====        srl s6, s7, ra
                                                  30'd    2357    : data = 32'h    7FDB80B7    ;    //    lui x1 523704      ====        lui ra, 523704
                                                  30'd    2358    : data = 32'h    01A7D733    ;    //    srl x14 x15 x26      ====        srl a4, a5, s10
                                                  30'd    2359    : data = 32'h    01D07933    ;    //    and x18 x0 x29      ====        and s2, zero, t4
                                                  30'd    2360    : data = 32'h    40550833    ;    //    sub x16 x10 x5      ====        sub a6, a0, t0
                                                  30'd    2361    : data = 32'h    33136E13    ;    //    ori x28 x6 817      ====        ori t3, t1, 817
                                                  30'd    2362    : data = 32'h    01ED9913    ;    //    slli x18 x27 30      ====        slli s2, s11, 30
                                                  30'd    2363    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2364    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2365    : data = 32'h    01F99193    ;    //    slli x3 x19 31      ====        slli gp, s3, 31
                                                  30'd    2366    : data = 32'h    015BC333    ;    //    xor x6 x23 x21      ====        xor t1, s7, s5
                                                  30'd    2367    : data = 32'h    6A506737    ;    //    lui x14 435462      ====        lui a4, 435462
                                                  30'd    2368    : data = 32'h    00B458B3    ;    //    srl x17 x8 x11      ====        srl a7, s0, a1
                                                  30'd    2369    : data = 32'h    94067597    ;    //    auipc x11 606311      ====        auipc a1, 606311
                                                  30'd    2370    : data = 32'h    6B190337    ;    //    lui x6 438672      ====        lui t1, 438672
                                                  30'd    2371    : data = 32'h    01DEDAB3    ;    //    srl x21 x29 x29      ====        srl s5, t4, t4
                                                  30'd    2372    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2373    : data = 32'h    00CF5A33    ;    //    srl x20 x30 x12      ====        srl s4, t5, a2
                                                  30'd    2374    : data = 32'h    A0EE8113    ;    //    addi x2 x29 -1522      ====        addi sp, t4, -1522
                                                  30'd    2375    : data = 32'h    00103CB3    ;    //    sltu x25 x0 x1      ====        sltu s9, zero, ra
                                                  30'd    2376    : data = 32'h    657F0C93    ;    //    addi x25 x30 1623      ====        addi s9, t5, 1623
                                                  30'd    2377    : data = 32'h    015F3AB3    ;    //    sltu x21 x30 x21      ====        sltu s5, t5, s5
                                                  30'd    2378    : data = 32'h    01D1FD33    ;    //    and x26 x3 x29      ====        and s10, gp, t4
                                                  30'd    2379    : data = 32'h    FB926893    ;    //    ori x17 x4 -71      ====        ori a7, tp, -71
                                                  30'd    2380    : data = 32'h    2563C793    ;    //    xori x15 x7 598      ====        xori a5, t2, 598
                                                  30'd    2381    : data = 32'h    CA322D37    ;    //    lui x26 828194      ====        lui s10, 828194
                                                  30'd    2382    : data = 32'h    00D08633    ;    //    add x12 x1 x13      ====        add a2, ra, a3
                                                  30'd    2383    : data = 32'h    B4B73093    ;    //    sltiu x1 x14 -1205      ====        sltiu ra, a4, -1205
                                                  30'd    2384    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2385    : data = 32'h    B3326D93    ;    //    ori x27 x4 -1229      ====        ori s11, tp, -1229
                                                  30'd    2386    : data = 32'h    521B3993    ;    //    sltiu x19 x22 1313      ====        sltiu s3, s6, 1313
                                                  30'd    2387    : data = 32'h    00C0FC33    ;    //    and x24 x1 x12      ====        and s8, ra, a2
                                                  30'd    2388    : data = 32'h    41F05933    ;    //    sra x18 x0 x31      ====        sra s2, zero, t6
                                                  30'd    2389    : data = 32'h    2DEB2013    ;    //    slti x0 x22 734      ====        slti zero, s6, 734
                                                  30'd    2390    : data = 32'h    012E9193    ;    //    slli x3 x29 18      ====        slli gp, t4, 18
                                                  30'd    2391    : data = 32'h    619D8A13    ;    //    addi x20 x27 1561      ====        addi s4, s11, 1561
                                                  30'd    2392    : data = 32'h    00C45E33    ;    //    srl x28 x8 x12      ====        srl t3, s0, a2
                                                  30'd    2393    : data = 32'h    95BF4BB7    ;    //    lui x23 613364      ====        lui s7, 613364
                                                  30'd    2394    : data = 32'h    0057D933    ;    //    srl x18 x15 x5      ====        srl s2, a5, t0
                                                  30'd    2395    : data = 32'h    DBD25C97    ;    //    auipc x25 900389      ====        auipc s9, 900389
                                                  30'd    2396    : data = 32'h    40C9DE33    ;    //    sra x28 x19 x12      ====        sra t3, s3, a2
                                                  30'd    2397    : data = 32'h    01A3D6B3    ;    //    srl x13 x7 x26      ====        srl a3, t2, s10
                                                  30'd    2398    : data = 32'h    62D60793    ;    //    addi x15 x12 1581      ====        addi a5, a2, 1581
                                                  30'd    2399    : data = 32'h    9EEF8EB7    ;    //    lui x29 651000      ====        lui t4, 651000
                                                  30'd    2400    : data = 32'h    01DED8B3    ;    //    srl x17 x29 x29      ====        srl a7, t4, t4
                                                  30'd    2401    : data = 32'h    01FABD33    ;    //    sltu x26 x21 x31      ====        sltu s10, s5, t6
                                                  30'd    2402    : data = 32'h    007E6433    ;    //    or x8 x28 x7      ====        or s0, t3, t2
                                                  30'd    2403    : data = 32'h    01D95E33    ;    //    srl x28 x18 x29      ====        srl t3, s2, t4
                                                  30'd    2404    : data = 32'h    406455B3    ;    //    sra x11 x8 x6      ====        sra a1, s0, t1
                                                  30'd    2405    : data = 32'h    B5E52A93    ;    //    slti x21 x10 -1186      ====        slti s5, a0, -1186
                                                  30'd    2406    : data = 32'h    01A717B3    ;    //    sll x15 x14 x26      ====        sll a5, a4, s10
                                                  30'd    2407    : data = 32'h    41B48833    ;    //    sub x16 x9 x27      ====        sub a6, s1, s11
                                                  30'd    2408    : data = 32'h    011E0133    ;    //    add x2 x28 x17      ====        add sp, t3, a7
                                                  30'd    2409    : data = 32'h    68663313    ;    //    sltiu x6 x12 1670      ====        sltiu t1, a2, 1670
                                                  30'd    2410    : data = 32'h    0003DD33    ;    //    srl x26 x7 x0      ====        srl s10, t2, zero
                                                  30'd    2411    : data = 32'h    E10C9DB7    ;    //    lui x27 921801      ====        lui s11, 921801
                                                  30'd    2412    : data = 32'h    223CF893    ;    //    andi x17 x25 547      ====        andi a7, s9, 547
                                                  30'd    2413    : data = 32'h    0152E0B3    ;    //    or x1 x5 x21      ====        or ra, t0, s5
                                                  30'd    2414    : data = 32'h    018A03B3    ;    //    add x7 x20 x24      ====        add t2, s4, s8
                                                  30'd    2415    : data = 32'h    40168D33    ;    //    sub x26 x13 x1      ====        sub s10, a3, ra
                                                  30'd    2416    : data = 32'h    09968C13    ;    //    addi x24 x13 153      ====        addi s8, a3, 153
                                                  30'd    2417    : data = 32'h    86AEAC93    ;    //    slti x25 x29 -1942      ====        slti s9, t4, -1942
                                                  30'd    2418    : data = 32'h    00E37A33    ;    //    and x20 x6 x14      ====        and s4, t1, a4
                                                  30'd    2419    : data = 32'h    81717613    ;    //    andi x12 x2 -2025      ====        andi a2, sp, -2025
                                                  30'd    2420    : data = 32'h    00F2C433    ;    //    xor x8 x5 x15      ====        xor s0, t0, a5
                                                  30'd    2421    : data = 32'h    01DAD333    ;    //    srl x6 x21 x29      ====        srl t1, s5, t4
                                                  30'd    2422    : data = 32'h    27342713    ;    //    slti x14 x8 627      ====        slti a4, s0, 627
                                                  30'd    2423    : data = 32'h    01CC1433    ;    //    sll x8 x24 x28      ====        sll s0, s8, t3
                                                  30'd    2424    : data = 32'h    BA6EE413    ;    //    ori x8 x29 -1114      ====        ori s0, t4, -1114
                                                  30'd    2425    : data = 32'h    015A55B3    ;    //    srl x11 x20 x21      ====        srl a1, s4, s5
                                                  30'd    2426    : data = 32'h    00486FB3    ;    //    or x31 x16 x4      ====        or t6, a6, tp
                                                  30'd    2427    : data = 32'h    833708B7    ;    //    lui x17 537456      ====        lui a7, 537456
                                                  30'd    2428    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2429    : data = 32'h    01861113    ;    //    slli x2 x12 24      ====        slli sp, a2, 24
                                                  30'd    2430    : data = 32'h    41A704B3    ;    //    sub x9 x14 x26      ====        sub s1, a4, s10
                                                  30'd    2431    : data = 32'h    0102AAB3    ;    //    slt x21 x5 x16      ====        slt s5, t0, a6
                                                  30'd    2432    : data = 32'h    019F5113    ;    //    srli x2 x30 25      ====        srli sp, t5, 25
                                                  30'd    2433    : data = 32'h    879B4A13    ;    //    xori x20 x22 -1927      ====        xori s4, s6, -1927
                                                  30'd    2434    : data = 32'h    147A7D13    ;    //    andi x26 x20 327      ====        andi s10, s4, 327
                                                  30'd    2435    : data = 32'h    258AB993    ;    //    sltiu x19 x21 600      ====        sltiu s3, s5, 600
                                                  30'd    2436    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2437    : data = 32'h    015317B3    ;    //    sll x15 x6 x21      ====        sll a5, t1, s5
                                                  30'd    2438    : data = 32'h    01643FB3    ;    //    sltu x31 x8 x22      ====        sltu t6, s0, s6
                                                  30'd    2439    : data = 32'h    014B65B3    ;    //    or x11 x22 x20      ====        or a1, s6, s4
                                                  30'd    2440    : data = 32'h    5A29F613    ;    //    andi x12 x19 1442      ====        andi a2, s3, 1442
                                                  30'd    2441    : data = 32'h    5863A413    ;    //    slti x8 x7 1414      ====        slti s0, t2, 1414
                                                  30'd    2442    : data = 32'h    30C3AB93    ;    //    slti x23 x7 780      ====        slti s7, t2, 780
                                                  30'd    2443    : data = 32'h    411DDA93    ;    //    srai x21 x27 17      ====        srai s5, s11, 17
                                                  30'd    2444    : data = 32'h    418FDE33    ;    //    sra x28 x31 x24      ====        sra t3, t6, s8
                                                  30'd    2445    : data = 32'h    FC2D4937    ;    //    lui x18 1032916      ====        lui s2, 1032916
                                                  30'd    2446    : data = 32'h    40AED793    ;    //    srai x15 x29 10      ====        srai a5, t4, 10
                                                  30'd    2447    : data = 32'h    25D2C793    ;    //    xori x15 x5 605      ====        xori a5, t0, 605
                                                  30'd    2448    : data = 32'h    6C20E937    ;    //    lui x18 442894      ====        lui s2, 442894
                                                  30'd    2449    : data = 32'h    F038B097    ;    //    auipc x1 983947      ====        auipc ra, 983947
                                                  30'd    2450    : data = 32'h    01B1DE13    ;    //    srli x28 x3 27      ====        srli t3, gp, 27
                                                  30'd    2451    : data = 32'h    3F150E17    ;    //    auipc x28 258384      ====        auipc t3, 258384
                                                  30'd    2452    : data = 32'h    A4FA6C13    ;    //    ori x24 x20 -1457      ====        ori s8, s4, -1457
                                                  30'd    2453    : data = 32'h    7C5D7193    ;    //    andi x3 x26 1989      ====        andi gp, s10, 1989
                                                  30'd    2454    : data = 32'h    0093D293    ;    //    srli x5 x7 9      ====        srli t0, t2, 9
                                                  30'd    2455    : data = 32'h    007CBE33    ;    //    sltu x28 x25 x7      ====        sltu t3, s9, t2
                                                  30'd    2456    : data = 32'h    7262C2B7    ;    //    lui x5 468524      ====        lui t0, 468524
                                                  30'd    2457    : data = 32'h    CE77E613    ;    //    ori x12 x15 -793      ====        ori a2, a5, -793
                                                  30'd    2458    : data = 32'h    00489AB3    ;    //    sll x21 x17 x4      ====        sll s5, a7, tp
                                                  30'd    2459    : data = 32'h    696BF813    ;    //    andi x16 x23 1686      ====        andi a6, s7, 1686
                                                  30'd    2460    : data = 32'h    CB086D93    ;    //    ori x27 x16 -848      ====        ori s11, a6, -848
                                                  30'd    2461    : data = 32'h    01AA9413    ;    //    slli x8 x21 26      ====        slli s0, s5, 26
                                                  30'd    2462    : data = 32'h    8EC84893    ;    //    xori x17 x16 -1812      ====        xori a7, a6, -1812
                                                  30'd    2463    : data = 32'h    0180F4B3    ;    //    and x9 x1 x24      ====        and s1, ra, s8
                                                  30'd    2464    : data = 32'h    00A309B3    ;    //    add x19 x6 x10      ====        add s3, t1, a0
                                                  30'd    2465    : data = 32'h    F52E4893    ;    //    xori x17 x28 -174      ====        xori a7, t3, -174
                                                  30'd    2466    : data = 32'h    012CB133    ;    //    sltu x2 x25 x18      ====        sltu sp, s9, s2
                                                  30'd    2467    : data = 32'h    02A1B293    ;    //    sltiu x5 x3 42      ====        sltiu t0, gp, 42
                                                  30'd    2468    : data = 32'h    15A7CFB7    ;    //    lui x31 88700      ====        lui t6, 88700
                                                  30'd    2469    : data = 32'h    00BEB813    ;    //    sltiu x16 x29 11      ====        sltiu a6, t4, 11
                                                  30'd    2470    : data = 32'h    401DD593    ;    //    srai x11 x27 1      ====        srai a1, s11, 1
                                                  30'd    2471    : data = 32'h    414CDFB3    ;    //    sra x31 x25 x20      ====        sra t6, s9, s4
                                                  30'd    2472    : data = 32'h    00EB1033    ;    //    sll x0 x22 x14      ====        sll zero, s6, a4
                                                  30'd    2473    : data = 32'h    7F9A6893    ;    //    ori x17 x20 2041      ====        ori a7, s4, 2041
                                                  30'd    2474    : data = 32'h    9EF7BD93    ;    //    sltiu x27 x15 -1553      ====        sltiu s11, a5, -1553
                                                  30'd    2475    : data = 32'h    01B99993    ;    //    slli x19 x19 27      ====        slli s3, s3, 27
                                                  30'd    2476    : data = 32'h    C6D97613    ;    //    andi x12 x18 -915      ====        andi a2, s2, -915
                                                  30'd    2477    : data = 32'h    01709E13    ;    //    slli x28 x1 23      ====        slli t3, ra, 23
                                                  30'd    2478    : data = 32'h    40B457B3    ;    //    sra x15 x8 x11      ====        sra a5, s0, a1
                                                  30'd    2479    : data = 32'h    001548B3    ;    //    xor x17 x10 x1      ====        xor a7, a0, ra
                                                  30'd    2480    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2481    : data = 32'h    00460DB3    ;    //    add x27 x12 x4      ====        add s11, a2, tp
                                                  30'd    2482    : data = 32'h    028C83B7    ;    //    lui x7 10440      ====        lui t2, 10440
                                                  30'd    2483    : data = 32'h    01BE03B3    ;    //    add x7 x28 x27      ====        add t2, t3, s11
                                                  30'd    2484    : data = 32'h    33708693    ;    //    addi x13 x1 823      ====        addi a3, ra, 823
                                                  30'd    2485    : data = 32'h    EA20AF93    ;    //    slti x31 x1 -350      ====        slti t6, ra, -350
                                                  30'd    2486    : data = 32'h    5F5B4D97    ;    //    auipc x27 390580      ====        auipc s11, 390580
                                                  30'd    2487    : data = 32'h    418B8333    ;    //    sub x6 x23 x24      ====        sub t1, s7, s8
                                                  30'd    2488    : data = 32'h    8D45C137    ;    //    lui x2 578652      ====        lui sp, 578652
                                                  30'd    2489    : data = 32'h    EE13A197    ;    //    auipc x3 975162      ====        auipc gp, 975162
                                                  30'd    2490    : data = 32'h    40FE81B3    ;    //    sub x3 x29 x15      ====        sub gp, t4, a5
                                                  30'd    2491    : data = 32'h    05F87A13    ;    //    andi x20 x16 95      ====        andi s4, a6, 95
                                                  30'd    2492    : data = 32'h    12B18D13    ;    //    addi x26 x3 299      ====        addi s10, gp, 299
                                                  30'd    2493    : data = 32'h    498B8E13    ;    //    addi x28 x23 1176      ====        addi t3, s7, 1176
                                                  30'd    2494    : data = 32'h    E356B113    ;    //    sltiu x2 x13 -459      ====        sltiu sp, a3, -459
                                                  30'd    2495    : data = 32'h    01B9ABB3    ;    //    slt x23 x19 x27      ====        slt s7, s3, s11
                                                  30'd    2496    : data = 32'h    7BCD6893    ;    //    ori x17 x26 1980      ====        ori a7, s10, 1980
                                                  30'd    2497    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2498    : data = 32'h    E90D7713    ;    //    andi x14 x26 -368      ====        andi a4, s10, -368
                                                  30'd    2499    : data = 32'h    06EC8193    ;    //    addi x3 x25 110      ====        addi gp, s9, 110
                                                  30'd    2500    : data = 32'h    017BCA33    ;    //    xor x20 x23 x23      ====        xor s4, s7, s7
                                                  30'd    2501    : data = 32'h    014E9193    ;    //    slli x3 x29 20      ====        slli gp, t4, 20
                                                  30'd    2502    : data = 32'h    4163D993    ;    //    srai x19 x7 22      ====        srai s3, t2, 22
                                                  30'd    2503    : data = 32'h    D35A0A93    ;    //    addi x21 x20 -715      ====        addi s5, s4, -715
                                                  30'd    2504    : data = 32'h    27AB3C97    ;    //    auipc x25 162483      ====        auipc s9, 162483
                                                  30'd    2505    : data = 32'h    E7D2C613    ;    //    xori x12 x5 -387      ====        xori a2, t0, -387
                                                  30'd    2506    : data = 32'h    01874133    ;    //    xor x2 x14 x24      ====        xor sp, a4, s8
                                                  30'd    2507    : data = 32'h    40715A33    ;    //    sra x20 x2 x7      ====        sra s4, sp, t2
                                                  30'd    2508    : data = 32'h    F4D5A313    ;    //    slti x6 x11 -179      ====        slti t1, a1, -179
                                                  30'd    2509    : data = 32'h    012C7BB3    ;    //    and x23 x24 x18      ====        and s7, s8, s2
                                                  30'd    2510    : data = 32'h    003E1FB3    ;    //    sll x31 x28 x3      ====        sll t6, t3, gp
                                                  30'd    2511    : data = 32'h    B3B2BE13    ;    //    sltiu x28 x5 -1221      ====        sltiu t3, t0, -1221
                                                  30'd    2512    : data = 32'h    01491833    ;    //    sll x16 x18 x20      ====        sll a6, s2, s4
                                                  30'd    2513    : data = 32'h    2396D117    ;    //    auipc x2 145773      ====        auipc sp, 145773
                                                  30'd    2514    : data = 32'h    41EA5333    ;    //    sra x6 x20 x30      ====        sra t1, s4, t5
                                                  30'd    2515    : data = 32'h    002BD6B3    ;    //    srl x13 x23 x2      ====        srl a3, s7, sp
                                                  30'd    2516    : data = 32'h    2C875097    ;    //    auipc x1 182389      ====        auipc ra, 182389
                                                  30'd    2517    : data = 32'h    0113C4B3    ;    //    xor x9 x7 x17      ====        xor s1, t2, a7
                                                  30'd    2518    : data = 32'h    C82FE313    ;    //    ori x6 x31 -894      ====        ori t1, t6, -894
                                                  30'd    2519    : data = 32'h    B8BBA697    ;    //    auipc x13 756666      ====        auipc a3, 756666
                                                  30'd    2520    : data = 32'h    00FEAAB3    ;    //    slt x21 x29 x15      ====        slt s5, t4, a5
                                                  30'd    2521    : data = 32'h    0153E1B3    ;    //    or x3 x7 x21      ====        or gp, t2, s5
                                                  30'd    2522    : data = 32'h    018B5033    ;    //    srl x0 x22 x24      ====        srl zero, s6, s8
                                                  30'd    2523    : data = 32'h    D0EFB193    ;    //    sltiu x3 x31 -754      ====        sltiu gp, t6, -754
                                                  30'd    2524    : data = 32'h    E2F30E13    ;    //    addi x28 x6 -465      ====        addi t3, t1, -465
                                                  30'd    2525    : data = 32'h    40F85333    ;    //    sra x6 x16 x15      ====        sra t1, a6, a5
                                                  30'd    2526    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2527    : data = 32'h    00ECE733    ;    //    or x14 x25 x14      ====        or a4, s9, a4
                                                  30'd    2528    : data = 32'h    01479413    ;    //    slli x8 x15 20      ====        slli s0, a5, 20
                                                  30'd    2529    : data = 32'h    00A2AE33    ;    //    slt x28 x5 x10      ====        slt t3, t0, a0
                                                  30'd    2530    : data = 32'h    38227B93    ;    //    andi x23 x4 898      ====        andi s7, tp, 898
                                                  30'd    2531    : data = 32'h    00505E33    ;    //    srl x28 x0 x5      ====        srl t3, zero, t0
                                                  30'd    2532    : data = 32'h    001D22B3    ;    //    slt x5 x26 x1      ====        slt t0, s10, ra
                                                  30'd    2533    : data = 32'h    0AF43093    ;    //    sltiu x1 x8 175      ====        sltiu ra, s0, 175
                                                  30'd    2534    : data = 32'h    00C1E333    ;    //    or x6 x3 x12      ====        or t1, gp, a2
                                                  30'd    2535    : data = 32'h    8626C593    ;    //    xori x11 x13 -1950      ====        xori a1, a3, -1950
                                                  30'd    2536    : data = 32'h    011D9113    ;    //    slli x2 x27 17      ====        slli sp, s11, 17
                                                  30'd    2537    : data = 32'h    CB504413    ;    //    xori x8 x0 -843      ====        xori s0, zero, -843
                                                  30'd    2538    : data = 32'h    89768093    ;    //    addi x1 x13 -1897      ====        addi ra, a3, -1897
                                                  30'd    2539    : data = 32'h    414C5C13    ;    //    srai x24 x24 20      ====        srai s8, s8, 20
                                                  30'd    2540    : data = 32'h    40CCDCB3    ;    //    sra x25 x25 x12      ====        sra s9, s9, a2
                                                  30'd    2541    : data = 32'h    B0520313    ;    //    addi x6 x4 -1275      ====        addi t1, tp, -1275
                                                  30'd    2542    : data = 32'h    004A9F93    ;    //    slli x31 x21 4      ====        slli t6, s5, 4
                                                  30'd    2543    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2544    : data = 32'h    40D95793    ;    //    srai x15 x18 13      ====        srai a5, s2, 13
                                                  30'd    2545    : data = 32'h    6A0B0E13    ;    //    addi x28 x22 1696      ====        addi t3, s6, 1696
                                                  30'd    2546    : data = 32'h    A9FAEC93    ;    //    ori x25 x21 -1377      ====        ori s9, s5, -1377
                                                  30'd    2547    : data = 32'h    AB337393    ;    //    andi x7 x6 -1357      ====        andi t2, t1, -1357
                                                  30'd    2548    : data = 32'h    016A9493    ;    //    slli x9 x21 22      ====        slli s1, s5, 22
                                                  30'd    2549    : data = 32'h    41670733    ;    //    sub x14 x14 x22      ====        sub a4, a4, s6
                                                  30'd    2550    : data = 32'h    004A3FB3    ;    //    sltu x31 x20 x4      ====        sltu t6, s4, tp
                                                  30'd    2551    : data = 32'h    01049033    ;    //    sll x0 x9 x16      ====        sll zero, s1, a6
                                                  30'd    2552    : data = 32'h    00E131B3    ;    //    sltu x3 x2 x14      ====        sltu gp, sp, a4
                                                  30'd    2553    : data = 32'h    00634CB3    ;    //    xor x25 x6 x6      ====        xor s9, t1, t1
                                                  30'd    2554    : data = 32'h    A9C74197    ;    //    auipc x3 695412      ====        auipc gp, 695412
                                                  30'd    2555    : data = 32'h    017F1813    ;    //    slli x16 x30 23      ====        slli a6, t5, 23
                                                  30'd    2556    : data = 32'h    E8E7FB13    ;    //    andi x22 x15 -370      ====        andi s6, a5, -370
                                                  30'd    2557    : data = 32'h    01F203B3    ;    //    add x7 x4 x31      ====        add t2, tp, t6
                                                  30'd    2558    : data = 32'h    010A94B3    ;    //    sll x9 x21 x16      ====        sll s1, s5, a6
                                                  30'd    2559    : data = 32'h    000CDF93    ;    //    srli x31 x25 0      ====        srli t6, s9, 0
                                                  30'd    2560    : data = 32'h    C3F37313    ;    //    andi x6 x6 -961      ====        andi t1, t1, -961
                                                  30'd    2561    : data = 32'h    CB428993    ;    //    addi x19 x5 -844      ====        addi s3, t0, -844
                                                  30'd    2562    : data = 32'h    236E3613    ;    //    sltiu x12 x28 566      ====        sltiu a2, t3, 566
                                                  30'd    2563    : data = 32'h    010E21B3    ;    //    slt x3 x28 x16      ====        slt gp, t3, a6
                                                  30'd    2564    : data = 32'h    C0EC4717    ;    //    auipc x14 790212      ====        auipc a4, 790212
                                                  30'd    2565    : data = 32'h    00799733    ;    //    sll x14 x19 x7      ====        sll a4, s3, t2
                                                  30'd    2566    : data = 32'h    00EC1193    ;    //    slli x3 x24 14      ====        slli gp, s8, 14
                                                  30'd    2567    : data = 32'h    01151593    ;    //    slli x11 x10 17      ====        slli a1, a0, 17
                                                  30'd    2568    : data = 32'h    CF0381B7    ;    //    lui x3 847928      ====        lui gp, 847928
                                                  30'd    2569    : data = 32'h    01685093    ;    //    srli x1 x16 22      ====        srli ra, a6, 22
                                                  30'd    2570    : data = 32'h    36130313    ;    //    addi x6 x6 865      ====        addi t1, t1, 865
                                                  30'd    2571    : data = 32'h    01A11BB3    ;    //    sll x23 x2 x26      ====        sll s7, sp, s10
                                                  30'd    2572    : data = 32'h    01799DB3    ;    //    sll x27 x19 x23      ====        sll s11, s3, s7
                                                  30'd    2573    : data = 32'h    B864A9B7    ;    //    lui x19 755274      ====        lui s3, 755274
                                                  30'd    2574    : data = 32'h    162D7413    ;    //    andi x8 x26 354      ====        andi s0, s10, 354
                                                  30'd    2575    : data = 32'h    594F0617    ;    //    auipc x12 365808      ====        auipc a2, 365808
                                                  30'd    2576    : data = 32'h    40F8D433    ;    //    sra x8 x17 x15      ====        sra s0, a7, a5
                                                  30'd    2577    : data = 32'h    01722CB3    ;    //    slt x25 x4 x23      ====        slt s9, tp, s7
                                                  30'd    2578    : data = 32'h    01255E13    ;    //    srli x28 x10 18      ====        srli t3, a0, 18
                                                  30'd    2579    : data = 32'h    69208F93    ;    //    addi x31 x1 1682      ====        addi t6, ra, 1682
                                                  30'd    2580    : data = 32'h    01E75D13    ;    //    srli x26 x14 30      ====        srli s10, a4, 30
                                                  30'd    2581    : data = 32'h    A51AF793    ;    //    andi x15 x21 -1455      ====        andi a5, s5, -1455
                                                  30'd    2582    : data = 32'h    017D7833    ;    //    and x16 x26 x23      ====        and a6, s10, s7
                                                  30'd    2583    : data = 32'h    A63D0837    ;    //    lui x16 680912      ====        lui a6, 680912
                                                  30'd    2584    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2585    : data = 32'h    84E2E413    ;    //    ori x8 x5 -1970      ====        ori s0, t0, -1970
                                                  30'd    2586    : data = 32'h    4104D137    ;    //    lui x2 266317      ====        lui sp, 266317
                                                  30'd    2587    : data = 32'h    5C67B913    ;    //    sltiu x18 x15 1478      ====        sltiu s2, a5, 1478
                                                  30'd    2588    : data = 32'h    D1A7BC37    ;    //    lui x24 858747      ====        li s8, 0xd1a7afde #start riscv_int_numeric_corner_stream_1
                                                  30'd    2589    : data = 32'h    FDEC0C13    ;    //    addi x24 x24 -34      ====        li s8, 0xd1a7afde #start riscv_int_numeric_corner_stream_1
                                                  30'd    2590    : data = 32'h    800003B7    ;    //    lui x7 524288      ====        li t2, 0x80000000
                                                  30'd    2591    : data = 32'h    00038393    ;    //    addi x7 x7 0      ====        li t2, 0x80000000
                                                  30'd    2592    : data = 32'h    800006B7    ;    //    lui x13 524288      ====        li a3, 0x80000000
                                                  30'd    2593    : data = 32'h    00068693    ;    //    addi x13 x13 0      ====        li a3, 0x80000000
                                                  30'd    2594    : data = 32'h    FFF00A13    ;    //    addi x20 x0 -1      ====        li s4, 0xffffffff
                                                  30'd    2595    : data = 32'h    00000913    ;    //    addi x18 x0 0      ====        li s2, 0x0
                                                  30'd    2596    : data = 32'h    FF9E0FB7    ;    //    lui x31 1047008      ====        li t6, 0xff9dfb64
                                                  30'd    2597    : data = 32'h    B64F8F93    ;    //    addi x31 x31 -1180      ====        li t6, 0xff9dfb64
                                                  30'd    2598    : data = 32'h    FFF00113    ;    //    addi x2 x0 -1      ====        li sp, 0xffffffff
                                                  30'd    2599    : data = 32'h    00000093    ;    //    addi x1 x0 0      ====        li ra, 0x0
                                                  30'd    2600    : data = 32'h    80000837    ;    //    lui x16 524288      ====        li a6, 0x80000000
                                                  30'd    2601    : data = 32'h    00080813    ;    //    addi x16 x16 0      ====        li a6, 0x80000000
                                                  30'd    2602    : data = 32'h    B2535E37    ;    //    lui x28 730421      ====        li t3, 0xb2534a0f
                                                  30'd    2603    : data = 32'h    A0FE0E13    ;    //    addi x28 x28 -1521      ====        li t3, 0xb2534a0f
                                                  30'd    2604    : data = 32'h    01F80E33    ;    //    add x28 x16 x31      ====        add t3, a6, t6
                                                  30'd    2605    : data = 32'h    041F8C13    ;    //    addi x24 x31 65      ====        addi s8, t6, 65
                                                  30'd    2606    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2607    : data = 32'h    7477B917    ;    //    auipc x18 477051      ====        auipc s2, 477051
                                                  30'd    2608    : data = 32'h    018E0C33    ;    //    add x24 x28 x24      ====        add s8, t3, s8
                                                  30'd    2609    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2610    : data = 32'h    01838933    ;    //    add x18 x7 x24      ====        add s2, t2, s8
                                                  30'd    2611    : data = 32'h    7B4956B7    ;    //    lui x13 504981      ====        lui a3, 504981
                                                  30'd    2612    : data = 32'h    002A0133    ;    //    add x2 x20 x2      ====        add sp, s4, sp
                                                  30'd    2613    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2614    : data = 32'h    40108E33    ;    //    sub x28 x1 x1      ====        sub t3, ra, ra
                                                  30'd    2615    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2616    : data = 32'h    00280FB3    ;    //    add x31 x16 x2      ====        add t6, a6, sp
                                                  30'd    2617    : data = 32'h    007A0E33    ;    //    add x28 x20 x7      ====        add t3, s4, t2
                                                  30'd    2618    : data = 32'h    EA4F8813    ;    //    addi x16 x31 -348      ====        addi a6, t6, -348
                                                  30'd    2619    : data = 32'h    002383B3    ;    //    add x7 x7 x2      ====        add t2, t2, sp
                                                  30'd    2620    : data = 32'h    1C008C13    ;    //    addi x24 x1 448      ====        addi s8, ra, 448
                                                  30'd    2621    : data = 32'h    FAB80113    ;    //    addi x2 x16 -85      ====        addi sp, a6, -85
                                                  30'd    2622    : data = 32'h    410803B3    ;    //    sub x7 x16 x16      ====        sub t2, a6, a6
                                                  30'd    2623    : data = 32'h    002C0FB3    ;    //    add x31 x24 x2      ====        add t6, s8, sp
                                                  30'd    2624    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2625    : data = 32'h    4D6E0093    ;    //    addi x1 x28 1238      ====        addi ra, t3, 1238
                                                  30'd    2626    : data = 32'h    402086B3    ;    //    sub x13 x1 x2      ====        sub a3, ra, sp
                                                  30'd    2627    : data = 32'h    410C00B3    ;    //    sub x1 x24 x16      ====        sub ra, s8, a6
                                                  30'd    2628    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2629    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2630    : data = 32'h    2B390813    ;    //    addi x16 x18 691      ====        addi a6, s2, 691
                                                  30'd    2631    : data = 32'h    401A0833    ;    //    sub x16 x20 x1      ====        sub a6, s4, ra
                                                  30'd    2632    : data = 32'h    F3DF0F97    ;    //    auipc x31 998896      ====        auipc t6, 998896
                                                  30'd    2633    : data = 32'h    5C5080EF    ;    //    jal x1 36292      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_1
                                                  30'd    2634    : data = 32'h    0039AFB3    ;    //    slt x31 x19 x3      ====        slt t6, s3, gp
                                                  30'd    2635    : data = 32'h    2C29C893    ;    //    xori x17 x19 706      ====        xori a7, s3, 706
                                                  30'd    2636    : data = 32'h    D5A1A397    ;    //    auipc x7 875034      ====        auipc t2, 875034
                                                  30'd    2637    : data = 32'h    00A759B3    ;    //    srl x19 x14 x10      ====        srl s3, a4, a0
                                                  30'd    2638    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2639    : data = 32'h    1AD2C293    ;    //    xori x5 x5 429      ====        xori t0, t0, 429
                                                  30'd    2640    : data = 32'h    40B85A33    ;    //    sra x20 x16 x11      ====        sra s4, a6, a1
                                                  30'd    2641    : data = 32'h    00DAE7B3    ;    //    or x15 x21 x13      ====        or a5, s5, a3
                                                  30'd    2642    : data = 32'h    877C5437    ;    //    lui x8 554949      ====        lui s0, 554949
                                                  30'd    2643    : data = 32'h    B4107D13    ;    //    andi x26 x0 -1215      ====        andi s10, zero, -1215
                                                  30'd    2644    : data = 32'h    00531633    ;    //    sll x12 x6 x5      ====        sll a2, t1, t0
                                                  30'd    2645    : data = 32'h    002FBD33    ;    //    sltu x26 x31 x2      ====        sltu s10, t6, sp
                                                  30'd    2646    : data = 32'h    007D6D33    ;    //    or x26 x26 x7      ====        or s10, s10, t2
                                                  30'd    2647    : data = 32'h    001EAFB3    ;    //    slt x31 x29 x1      ====        slt t6, t4, ra
                                                  30'd    2648    : data = 32'h    0DD97C93    ;    //    andi x25 x18 221      ====        andi s9, s2, 221
                                                  30'd    2649    : data = 32'h    408DD293    ;    //    srai x5 x27 8      ====        srai t0, s11, 8
                                                  30'd    2650    : data = 32'h    40D0D733    ;    //    sra x14 x1 x13      ====        sra a4, ra, a3
                                                  30'd    2651    : data = 32'h    016FF8B3    ;    //    and x17 x31 x22      ====        and a7, t6, s6
                                                  30'd    2652    : data = 32'h    01CD6633    ;    //    or x12 x26 x28      ====        or a2, s10, t3
                                                  30'd    2653    : data = 32'h    842DE913    ;    //    ori x18 x27 -1982      ====        ori s2, s11, -1982
                                                  30'd    2654    : data = 32'h    4107D2B3    ;    //    sra x5 x15 x16      ====        sra t0, a5, a6
                                                  30'd    2655    : data = 32'h    9EE08E93    ;    //    addi x29 x1 -1554      ====        addi t4, ra, -1554
                                                  30'd    2656    : data = 32'h    01B095B3    ;    //    sll x11 x1 x27      ====        sll a1, ra, s11
                                                  30'd    2657    : data = 32'h    008B6DB3    ;    //    or x27 x22 x8      ====        or s11, s6, s0
                                                  30'd    2658    : data = 32'h    00E59333    ;    //    sll x6 x11 x14      ====        sll t1, a1, a4
                                                  30'd    2659    : data = 32'h    00DFD013    ;    //    srli x0 x31 13      ====        srli zero, t6, 13
                                                  30'd    2660    : data = 32'h    01574A33    ;    //    xor x20 x14 x21      ====        xor s4, a4, s5
                                                  30'd    2661    : data = 32'h    40D35133    ;    //    sra x2 x6 x13      ====        sra sp, t1, a3
                                                  30'd    2662    : data = 32'h    000BB933    ;    //    sltu x18 x23 x0      ====        sltu s2, s7, zero
                                                  30'd    2663    : data = 32'h    A4DCC013    ;    //    xori x0 x25 -1459      ====        xori zero, s9, -1459
                                                  30'd    2664    : data = 32'h    018AD593    ;    //    srli x11 x21 24      ====        srli a1, s5, 24
                                                  30'd    2665    : data = 32'h    B33EC493    ;    //    xori x9 x29 -1229      ====        xori s1, t4, -1229
                                                  30'd    2666    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2667    : data = 32'h    001F1EB3    ;    //    sll x29 x30 x1      ====        sll t4, t5, ra
                                                  30'd    2668    : data = 32'h    012B5833    ;    //    srl x16 x22 x18      ====        srl a6, s6, s2
                                                  30'd    2669    : data = 32'h    01E37A33    ;    //    and x20 x6 x30      ====        and s4, t1, t5
                                                  30'd    2670    : data = 32'h    7C8EC113    ;    //    xori x2 x29 1992      ====        xori sp, t4, 1992
                                                  30'd    2671    : data = 32'h    00A69933    ;    //    sll x18 x13 x10      ====        sll s2, a3, a0
                                                  30'd    2672    : data = 32'h    3F437A93    ;    //    andi x21 x6 1012      ====        andi s5, t1, 1012
                                                  30'd    2673    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2674    : data = 32'h    D76AF897    ;    //    auipc x17 882351      ====        auipc a7, 882351
                                                  30'd    2675    : data = 32'h    01994B33    ;    //    xor x22 x18 x25      ====        xor s6, s2, s9
                                                  30'd    2676    : data = 32'h    37616313    ;    //    ori x6 x2 886      ====        ori t1, sp, 886
                                                  30'd    2677    : data = 32'h    40298EB3    ;    //    sub x29 x19 x2      ====        sub t4, s3, sp
                                                  30'd    2678    : data = 32'h    415AD1B3    ;    //    sra x3 x21 x21      ====        sra gp, s5, s5
                                                  30'd    2679    : data = 32'h    000477B3    ;    //    and x15 x8 x0      ====        and a5, s0, zero
                                                  30'd    2680    : data = 32'h    CAB0F813    ;    //    andi x16 x1 -853      ====        andi a6, ra, -853
                                                  30'd    2681    : data = 32'h    004D6333    ;    //    or x6 x26 x4      ====        or t1, s10, tp
                                                  30'd    2682    : data = 32'h    5ACA3693    ;    //    sltiu x13 x20 1452      ====        sltiu a3, s4, 1452
                                                  30'd    2683    : data = 32'h    0143B733    ;    //    sltu x14 x7 x20      ====        sltu a4, t2, s4
                                                  30'd    2684    : data = 32'h    1A524313    ;    //    xori x6 x4 421      ====        xori t1, tp, 421
                                                  30'd    2685    : data = 32'h    00EA9C13    ;    //    slli x24 x21 14      ====        slli s8, s5, 14
                                                  30'd    2686    : data = 32'h    222ECA93    ;    //    xori x21 x29 546      ====        xori s5, t4, 546
                                                  30'd    2687    : data = 32'h    41915E33    ;    //    sra x28 x2 x25      ====        sra t3, sp, s9
                                                  30'd    2688    : data = 32'h    6478EB13    ;    //    ori x22 x17 1607      ====        ori s6, a7, 1607
                                                  30'd    2689    : data = 32'h    E4C56A13    ;    //    ori x20 x10 -436      ====        ori s4, a0, -436
                                                  30'd    2690    : data = 32'h    01AB5D33    ;    //    srl x26 x22 x26      ====        srl s10, s6, s10
                                                  30'd    2691    : data = 32'h    8953A293    ;    //    slti x5 x7 -1899      ====        slti t0, t2, -1899
                                                  30'd    2692    : data = 32'h    415A0933    ;    //    sub x18 x20 x21      ====        sub s2, s4, s5
                                                  30'd    2693    : data = 32'h    0542A2B7    ;    //    lui x5 21546      ====        lui t0, 21546
                                                  30'd    2694    : data = 32'h    011015B3    ;    //    sll x11 x0 x17      ====        sll a1, zero, a7
                                                  30'd    2695    : data = 32'h    00929993    ;    //    slli x19 x5 9      ====        slli s3, t0, 9
                                                  30'd    2696    : data = 32'h    407AD493    ;    //    srai x9 x21 7      ====        srai s1, s5, 7
                                                  30'd    2697    : data = 32'h    00DA5CB3    ;    //    srl x25 x20 x13      ====        srl s9, s4, a3
                                                  30'd    2698    : data = 32'h    261B8F93    ;    //    addi x31 x23 609      ====        addi t6, s7, 609
                                                  30'd    2699    : data = 32'h    FAE10413    ;    //    addi x8 x2 -82      ====        addi s0, sp, -82
                                                  30'd    2700    : data = 32'h    01907AB3    ;    //    and x21 x0 x25      ====        and s5, zero, s9
                                                  30'd    2701    : data = 32'h    01A03933    ;    //    sltu x18 x0 x26      ====        sltu s2, zero, s10
                                                  30'd    2702    : data = 32'h    9A578913    ;    //    addi x18 x15 -1627      ====        addi s2, a5, -1627
                                                  30'd    2703    : data = 32'h    0033ABB3    ;    //    slt x23 x7 x3      ====        slt s7, t2, gp
                                                  30'd    2704    : data = 32'h    01702EB3    ;    //    slt x29 x0 x23      ====        slt t4, zero, s7
                                                  30'd    2705    : data = 32'h    53BCBD13    ;    //    sltiu x26 x25 1339      ====        sltiu s10, s9, 1339
                                                  30'd    2706    : data = 32'h    00711033    ;    //    sll x0 x2 x7      ====        sll zero, sp, t2
                                                  30'd    2707    : data = 32'h    01966633    ;    //    or x12 x12 x25      ====        or a2, a2, s9
                                                  30'd    2708    : data = 32'h    40305813    ;    //    srai x16 x0 3      ====        srai a6, zero, 3
                                                  30'd    2709    : data = 32'h    E4AC6D13    ;    //    ori x26 x24 -438      ====        ori s10, s8, -438
                                                  30'd    2710    : data = 32'h    01399413    ;    //    slli x8 x19 19      ====        slli s0, s3, 19
                                                  30'd    2711    : data = 32'h    9109EB13    ;    //    ori x22 x19 -1776      ====        ori s6, s3, -1776
                                                  30'd    2712    : data = 32'h    ABA7BA97    ;    //    auipc x21 703099      ====        auipc s5, 703099
                                                  30'd    2713    : data = 32'h    011DD1B3    ;    //    srl x3 x27 x17      ====        srl gp, s11, a7
                                                  30'd    2714    : data = 32'h    011F9CB3    ;    //    sll x25 x31 x17      ====        sll s9, t6, a7
                                                  30'd    2715    : data = 32'h    01EAF333    ;    //    and x6 x21 x30      ====        and t1, s5, t5
                                                  30'd    2716    : data = 32'h    010D9133    ;    //    sll x2 x27 x16      ====        sll sp, s11, a6
                                                  30'd    2717    : data = 32'h    83D5ED93    ;    //    ori x27 x11 -1987      ====        ori s11, a1, -1987
                                                  30'd    2718    : data = 32'h    A71CE293    ;    //    ori x5 x25 -1423      ====        ori t0, s9, -1423
                                                  30'd    2719    : data = 32'h    00401913    ;    //    slli x18 x0 4      ====        slli s2, zero, 4
                                                  30'd    2720    : data = 32'h    01A31713    ;    //    slli x14 x6 26      ====        slli a4, t1, 26
                                                  30'd    2721    : data = 32'h    014B4333    ;    //    xor x6 x22 x20      ====        xor t1, s6, s4
                                                  30'd    2722    : data = 32'h    005F5C13    ;    //    srli x24 x30 5      ====        srli s8, t5, 5
                                                  30'd    2723    : data = 32'h    01092B37    ;    //    lui x22 4242      ====        lui s6, 4242
                                                  30'd    2724    : data = 32'h    401456B3    ;    //    sra x13 x8 x1      ====        sra a3, s0, ra
                                                  30'd    2725    : data = 32'h    00EF44B3    ;    //    xor x9 x30 x14      ====        xor s1, t5, a4
                                                  30'd    2726    : data = 32'h    41BFDC33    ;    //    sra x24 x31 x27      ====        sra s8, t6, s11
                                                  30'd    2727    : data = 32'h    01C219B3    ;    //    sll x19 x4 x28      ====        sll s3, tp, t3
                                                  30'd    2728    : data = 32'h    BB5BFD17    ;    //    auipc x26 767423      ====        auipc s10, 767423
                                                  30'd    2729    : data = 32'h    01A3D433    ;    //    srl x8 x7 x26      ====        srl s0, t2, s10
                                                  30'd    2730    : data = 32'h    011AB133    ;    //    sltu x2 x21 x17      ====        sltu sp, s5, a7
                                                  30'd    2731    : data = 32'h    DA3B8C13    ;    //    addi x24 x23 -605      ====        addi s8, s7, -605
                                                  30'd    2732    : data = 32'h    018F60B3    ;    //    or x1 x30 x24      ====        or ra, t5, s8
                                                  30'd    2733    : data = 32'h    A3D115B7    ;    //    lui x11 670993      ====        lui a1, 670993
                                                  30'd    2734    : data = 32'h    4C094C13    ;    //    xori x24 x18 1216      ====        xori s8, s2, 1216
                                                  30'd    2735    : data = 32'h    74A6E193    ;    //    ori x3 x13 1866      ====        ori gp, a3, 1866
                                                  30'd    2736    : data = 32'h    019A20B3    ;    //    slt x1 x20 x25      ====        slt ra, s4, s9
                                                  30'd    2737    : data = 32'h    00E49193    ;    //    slli x3 x9 14      ====        slli gp, s1, 14
                                                  30'd    2738    : data = 32'h    005085B3    ;    //    add x11 x1 x5      ====        add a1, ra, t0
                                                  30'd    2739    : data = 32'h    B7A7C613    ;    //    xori x12 x15 -1158      ====        xori a2, a5, -1158
                                                  30'd    2740    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2741    : data = 32'h    F63D1F97    ;    //    auipc x31 1008593      ====        auipc t6, 1008593
                                                  30'd    2742    : data = 32'h    0E5FFB93    ;    //    andi x23 x31 229      ====        andi s7, t6, 229
                                                  30'd    2743    : data = 32'h    40095093    ;    //    srai x1 x18 0      ====        srai ra, s2, 0
                                                  30'd    2744    : data = 32'h    00FDDD13    ;    //    srli x26 x27 15      ====        srli s10, s11, 15
                                                  30'd    2745    : data = 32'h    7F0E6693    ;    //    ori x13 x28 2032      ====        ori a3, t3, 2032
                                                  30'd    2746    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2747    : data = 32'h    89FA3713    ;    //    sltiu x14 x20 -1889      ====        sltiu a4, s4, -1889
                                                  30'd    2748    : data = 32'h    14EA0A93    ;    //    addi x21 x20 334      ====        addi s5, s4, 334
                                                  30'd    2749    : data = 32'h    01D13093    ;    //    sltiu x1 x2 29      ====        sltiu ra, sp, 29
                                                  30'd    2750    : data = 32'h    0402F013    ;    //    andi x0 x5 64      ====        andi zero, t0, 64
                                                  30'd    2751    : data = 32'h    36E26937    ;    //    lui x18 224806      ====        lui s2, 224806
                                                  30'd    2752    : data = 32'h    01803633    ;    //    sltu x12 x0 x24      ====        sltu a2, zero, s8
                                                  30'd    2753    : data = 32'h    5D86E1B7    ;    //    lui x3 383086      ====        lui gp, 383086
                                                  30'd    2754    : data = 32'h    E15E2713    ;    //    slti x14 x28 -491      ====        slti a4, t3, -491
                                                  30'd    2755    : data = 32'h    401755B3    ;    //    sra x11 x14 x1      ====        sra a1, a4, ra
                                                  30'd    2756    : data = 32'h    411153B3    ;    //    sra x7 x2 x17      ====        sra t2, sp, a7
                                                  30'd    2757    : data = 32'h    096B7813    ;    //    andi x16 x22 150      ====        andi a6, s6, 150
                                                  30'd    2758    : data = 32'h    0106E133    ;    //    or x2 x13 x16      ====        or sp, a3, a6
                                                  30'd    2759    : data = 32'h    417E0DB3    ;    //    sub x27 x28 x23      ====        sub s11, t3, s7
                                                  30'd    2760    : data = 32'h    01F41D33    ;    //    sll x26 x8 x31      ====        sll s10, s0, t6
                                                  30'd    2761    : data = 32'h    0045D293    ;    //    srli x5 x11 4      ====        srli t0, a1, 4
                                                  30'd    2762    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2763    : data = 32'h    013CA0B3    ;    //    slt x1 x25 x19      ====        slt ra, s9, s3
                                                  30'd    2764    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2765    : data = 32'h    0150CFB3    ;    //    xor x31 x1 x21      ====        xor t6, ra, s5
                                                  30'd    2766    : data = 32'h    5B24EC13    ;    //    ori x24 x9 1458      ====        ori s8, s1, 1458
                                                  30'd    2767    : data = 32'h    01EB9113    ;    //    slli x2 x23 30      ====        slli sp, s7, 30
                                                  30'd    2768    : data = 32'h    211AC293    ;    //    xori x5 x21 529      ====        xori t0, s5, 529
                                                  30'd    2769    : data = 32'h    0100F5B3    ;    //    and x11 x1 x16      ====        and a1, ra, a6
                                                  30'd    2770    : data = 32'h    4126D813    ;    //    srai x16 x13 18      ====        srai a6, a3, 18
                                                  30'd    2771    : data = 32'h    02E20817    ;    //    auipc x16 11808      ====        auipc a6, 11808
                                                  30'd    2772    : data = 32'h    406C5393    ;    //    srai x7 x24 6      ====        srai t2, s8, 6
                                                  30'd    2773    : data = 32'h    40BA0733    ;    //    sub x14 x20 x11      ====        sub a4, s4, a1
                                                  30'd    2774    : data = 32'h    408A5F93    ;    //    srai x31 x20 8      ====        srai t6, s4, 8
                                                  30'd    2775    : data = 32'h    6689B817    ;    //    auipc x16 419995      ====        auipc a6, 419995
                                                  30'd    2776    : data = 32'h    00EEECB3    ;    //    or x25 x29 x14      ====        or s9, t4, a4
                                                  30'd    2777    : data = 32'h    7C480D13    ;    //    addi x26 x16 1988      ====        addi s10, a6, 1988
                                                  30'd    2778    : data = 32'h    41EDD6B3    ;    //    sra x13 x27 x30      ====        sra a3, s11, t5
                                                  30'd    2779    : data = 32'h    00F26133    ;    //    or x2 x4 x15      ====        or sp, tp, a5
                                                  30'd    2780    : data = 32'h    01C37733    ;    //    and x14 x6 x28      ====        and a4, t1, t3
                                                  30'd    2781    : data = 32'h    00B164B3    ;    //    or x9 x2 x11      ====        or s1, sp, a1
                                                  30'd    2782    : data = 32'h    00F37833    ;    //    and x16 x6 x15      ====        and a6, t1, a5
                                                  30'd    2783    : data = 32'h    139EE313    ;    //    ori x6 x29 313      ====        ori t1, t4, 313
                                                  30'd    2784    : data = 32'h    010C5593    ;    //    srli x11 x24 16      ====        srli a1, s8, 16
                                                  30'd    2785    : data = 32'h    009B80B3    ;    //    add x1 x23 x9      ====        add ra, s7, s1
                                                  30'd    2786    : data = 32'h    01EFCFB3    ;    //    xor x31 x31 x30      ====        xor t6, t6, t5
                                                  30'd    2787    : data = 32'h    B128F193    ;    //    andi x3 x17 -1262      ====        andi gp, a7, -1262
                                                  30'd    2788    : data = 32'h    00DD5993    ;    //    srli x19 x26 13      ====        srli s3, s10, 13
                                                  30'd    2789    : data = 32'h    01CF12B3    ;    //    sll x5 x30 x28      ====        sll t0, t5, t3
                                                  30'd    2790    : data = 32'h    D894C293    ;    //    xori x5 x9 -631      ====        xori t0, s1, -631
                                                  30'd    2791    : data = 32'h    40F15AB3    ;    //    sra x21 x2 x15      ====        sra s5, sp, a5
                                                  30'd    2792    : data = 32'h    00360A33    ;    //    add x20 x12 x3      ====        add s4, a2, gp
                                                  30'd    2793    : data = 32'h    D3136713    ;    //    ori x14 x6 -719      ====        ori a4, t1, -719
                                                  30'd    2794    : data = 32'h    01DF6433    ;    //    or x8 x30 x29      ====        or s0, t5, t4
                                                  30'd    2795    : data = 32'h    155EF313    ;    //    andi x6 x29 341      ====        andi t1, t4, 341
                                                  30'd    2796    : data = 32'h    015C53B3    ;    //    srl x7 x24 x21      ====        srl t2, s8, s5
                                                  30'd    2797    : data = 32'h    524C6E93    ;    //    ori x29 x24 1316      ====        ori t4, s8, 1316
                                                  30'd    2798    : data = 32'h    00C3C1B3    ;    //    xor x3 x7 x12      ====        xor gp, t2, a2
                                                  30'd    2799    : data = 32'h    40CBD713    ;    //    srai x14 x23 12      ====        srai a4, s7, 12
                                                  30'd    2800    : data = 32'h    00E6EA93    ;    //    ori x21 x13 14      ====        ori s5, a3, 14
                                                  30'd    2801    : data = 32'h    BC232293    ;    //    slti x5 x6 -1086      ====        slti t0, t1, -1086
                                                  30'd    2802    : data = 32'h    01C9DA13    ;    //    srli x20 x19 28      ====        srli s4, s3, 28
                                                  30'd    2803    : data = 32'h    00B78833    ;    //    add x16 x15 x11      ====        add a6, a5, a1
                                                  30'd    2804    : data = 32'h    019D5FB3    ;    //    srl x31 x26 x25      ====        srl t6, s10, s9
                                                  30'd    2805    : data = 32'h    60E3AA13    ;    //    slti x20 x7 1550      ====        slti s4, t2, 1550
                                                  30'd    2806    : data = 32'h    FE0EFF93    ;    //    andi x31 x29 -32      ====        andi t6, t4, -32
                                                  30'd    2807    : data = 32'h    005DDC13    ;    //    srli x24 x27 5      ====        srli s8, s11, 5
                                                  30'd    2808    : data = 32'h    3BD92293    ;    //    slti x5 x18 957      ====        slti t0, s2, 957
                                                  30'd    2809    : data = 32'h    FFF00A13    ;    //    addi x20 x0 -1      ====        li s4, 0xffffffff #start riscv_int_numeric_corner_stream_16
                                                  30'd    2810    : data = 32'h    48D052B7    ;    //    lui x5 298245      ====        li t0, 0x48d05214
                                                  30'd    2811    : data = 32'h    21428293    ;    //    addi x5 x5 532      ====        li t0, 0x48d05214
                                                  30'd    2812    : data = 32'h    800001B7    ;    //    lui x3 524288      ====        li gp, 0x80000000
                                                  30'd    2813    : data = 32'h    00018193    ;    //    addi x3 x3 0      ====        li gp, 0x80000000
                                                  30'd    2814    : data = 32'h    639FCBB7    ;    //    lui x23 408060      ====        li s7, 0x639fc7a7
                                                  30'd    2815    : data = 32'h    7A7B8B93    ;    //    addi x23 x23 1959      ====        li s7, 0x639fc7a7
                                                  30'd    2816    : data = 32'h    00000613    ;    //    addi x12 x0 0      ====        li a2, 0x0
                                                  30'd    2817    : data = 32'h    80000137    ;    //    lui x2 524288      ====        li sp, 0x80000000
                                                  30'd    2818    : data = 32'h    00010113    ;    //    addi x2 x2 0      ====        li sp, 0x80000000
                                                  30'd    2819    : data = 32'h    F036A437    ;    //    lui x8 983914      ====        li s0, 0xf036a43d
                                                  30'd    2820    : data = 32'h    43D40413    ;    //    addi x8 x8 1085      ====        li s0, 0xf036a43d
                                                  30'd    2821    : data = 32'h    500777B7    ;    //    lui x15 327799      ====        li a5, 0x5007745e
                                                  30'd    2822    : data = 32'h    45E78793    ;    //    addi x15 x15 1118      ====        li a5, 0x5007745e
                                                  30'd    2823    : data = 32'h    FFF00493    ;    //    addi x9 x0 -1      ====        li s1, 0xffffffff
                                                  30'd    2824    : data = 32'h    BCF35C37    ;    //    lui x24 773941      ====        li s8, 0xbcf34c4c
                                                  30'd    2825    : data = 32'h    C4CC0C13    ;    //    addi x24 x24 -948      ====        li s8, 0xbcf34c4c
                                                  30'd    2826    : data = 32'h    40310133    ;    //    sub x2 x2 x3      ====        sub sp, sp, gp
                                                  30'd    2827    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2828    : data = 32'h    D5C614B7    ;    //    lui x9 875617      ====        lui s1, 875617
                                                  30'd    2829    : data = 32'h    018782B3    ;    //    add x5 x15 x24      ====        add t0, a5, s8
                                                  30'd    2830    : data = 32'h    417B8BB3    ;    //    sub x23 x23 x23      ====        sub s7, s7, s7
                                                  30'd    2831    : data = 32'h    9B827117    ;    //    auipc x2 636967      ====        auipc sp, 636967
                                                  30'd    2832    : data = 32'h    FEA75C37    ;    //    lui x24 1043061      ====        lui s8, 1043061
                                                  30'd    2833    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2834    : data = 32'h    40F18BB3    ;    //    sub x23 x3 x15      ====        sub s7, gp, a5
                                                  30'd    2835    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2836    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2837    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2838    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2839    : data = 32'h    418A07B3    ;    //    sub x15 x20 x24      ====        sub a5, s4, s8
                                                  30'd    2840    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2841    : data = 32'h    00948A33    ;    //    add x20 x9 x9      ====        add s4, s1, s1
                                                  30'd    2842    : data = 32'h    40310C33    ;    //    sub x24 x2 x3      ====        sub s8, sp, gp
                                                  30'd    2843    : data = 32'h    9B240493    ;    //    addi x9 x8 -1614      ====        addi s1, s0, -1614
                                                  30'd    2844    : data = 32'h    5DF09197    ;    //    auipc x3 384777      ====        auipc gp, 384777
                                                  30'd    2845    : data = 32'h    16DFABB7    ;    //    lui x23 93690      ====        lui s7, 93690
                                                  30'd    2846    : data = 32'h    D58A0A13    ;    //    addi x20 x20 -680      ====        addi s4, s4, -680
                                                  30'd    2847    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2848    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2849    : data = 32'h    5A979497    ;    //    auipc x9 371065      ====        auipc s1, 371065
                                                  30'd    2850    : data = 32'h    36848C13    ;    //    addi x24 x9 872      ====        addi s8, s1, 872
                                                  30'd    2851    : data = 32'h    01848A33    ;    //    add x20 x9 x24      ====        add s4, s1, s8
                                                  30'd    2852    : data = 32'h    6E8924B7    ;    //    lui x9 452754      ====        lui s1, 452754
                                                  30'd    2853    : data = 32'h    F37A0413    ;    //    addi x8 x20 -201      ====        addi s0, s4, -201
                                                  30'd    2854    : data = 32'h    018104B3    ;    //    add x9 x2 x24      ====        add s1, sp, s8
                                                  30'd    2855    : data = 32'h    417182B3    ;    //    sub x5 x3 x23      ====        sub t0, gp, s7
                                                  30'd    2856    : data = 32'h    249080EF    ;    //    jal x1 35400      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_16
                                                  30'd    2857    : data = 32'h    415E5A13    ;    //    srai x20 x28 21      ====        srai s4, t3, 21
                                                  30'd    2858    : data = 32'h    01299CB3    ;    //    sll x25 x19 x18      ====        sll s9, s3, s2
                                                  30'd    2859    : data = 32'h    017FC2B3    ;    //    xor x5 x31 x23      ====        xor t0, t6, s7
                                                  30'd    2860    : data = 32'h    0FDCE093    ;    //    ori x1 x25 253      ====        ori ra, s9, 253
                                                  30'd    2861    : data = 32'h    B2284013    ;    //    xori x0 x16 -1246      ====        xori zero, a6, -1246
                                                  30'd    2862    : data = 32'h    00CA1913    ;    //    slli x18 x20 12      ====        slli s2, s4, 12
                                                  30'd    2863    : data = 32'h    3D0A7B13    ;    //    andi x22 x20 976      ====        andi s6, s4, 976
                                                  30'd    2864    : data = 32'h    6CF23393    ;    //    sltiu x7 x4 1743      ====        sltiu t2, tp, 1743
                                                  30'd    2865    : data = 32'h    56127793    ;    //    andi x15 x4 1377      ====        andi a5, tp, 1377
                                                  30'd    2866    : data = 32'h    00CB29B3    ;    //    slt x19 x22 x12      ====        slt s3, s6, a2
                                                  30'd    2867    : data = 32'h    00007AB3    ;    //    and x21 x0 x0      ====        and s5, zero, zero
                                                  30'd    2868    : data = 32'h    01BF8A33    ;    //    add x20 x31 x27      ====        add s4, t6, s11
                                                  30'd    2869    : data = 32'h    426ABB17    ;    //    auipc x22 272043      ====        auipc s6, 272043
                                                  30'd    2870    : data = 32'h    D3363C13    ;    //    sltiu x24 x12 -717      ====        sltiu s8, a2, -717
                                                  30'd    2871    : data = 32'h    00815AB3    ;    //    srl x21 x2 x8      ====        srl s5, sp, s0
                                                  30'd    2872    : data = 32'h    C9BF4693    ;    //    xori x13 x30 -869      ====        xori a3, t5, -869
                                                  30'd    2873    : data = 32'h    3597F713    ;    //    andi x14 x15 857      ====        andi a4, a5, 857
                                                  30'd    2874    : data = 32'h    00999793    ;    //    slli x15 x19 9      ====        slli a5, s3, 9
                                                  30'd    2875    : data = 32'h    00D75F93    ;    //    srli x31 x14 13      ====        srli t6, a4, 13
                                                  30'd    2876    : data = 32'h    00036BB3    ;    //    or x23 x6 x0      ====        or s7, t1, zero
                                                  30'd    2877    : data = 32'h    002A6CB3    ;    //    or x25 x20 x2      ====        or s9, s4, sp
                                                  30'd    2878    : data = 32'h    01F95D93    ;    //    srli x27 x18 31      ====        srli s11, s2, 31
                                                  30'd    2879    : data = 32'h    01CCEB33    ;    //    or x22 x25 x28      ====        or s6, s9, t3
                                                  30'd    2880    : data = 32'h    4EECBF93    ;    //    sltiu x31 x25 1262      ====        sltiu t6, s9, 1262
                                                  30'd    2881    : data = 32'h    C28D8A13    ;    //    addi x20 x27 -984      ====        addi s4, s11, -984
                                                  30'd    2882    : data = 32'h    40EB83B3    ;    //    sub x7 x23 x14      ====        sub t2, s7, a4
                                                  30'd    2883    : data = 32'h    412D00B3    ;    //    sub x1 x26 x18      ====        sub ra, s10, s2
                                                  30'd    2884    : data = 32'h    00AE80B3    ;    //    add x1 x29 x10      ====        add ra, t4, a0
                                                  30'd    2885    : data = 32'h    00BDD033    ;    //    srl x0 x27 x11      ====        srl zero, s11, a1
                                                  30'd    2886    : data = 32'h    01A91593    ;    //    slli x11 x18 26      ====        slli a1, s2, 26
                                                  30'd    2887    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2888    : data = 32'h    41325F93    ;    //    srai x31 x4 19      ====        srai t6, tp, 19
                                                  30'd    2889    : data = 32'h    00140333    ;    //    add x6 x8 x1      ====        add t1, s0, ra
                                                  30'd    2890    : data = 32'h    11D3F193    ;    //    andi x3 x7 285      ====        andi gp, t2, 285
                                                  30'd    2891    : data = 32'h    0053FAB3    ;    //    and x21 x7 x5      ====        and s5, t2, t0
                                                  30'd    2892    : data = 32'h    98283713    ;    //    sltiu x14 x16 -1662      ====        sltiu a4, a6, -1662
                                                  30'd    2893    : data = 32'h    410CD993    ;    //    srai x19 x25 16      ====        srai s3, s9, 16
                                                  30'd    2894    : data = 32'h    0011D793    ;    //    srli x15 x3 1      ====        srli a5, gp, 1
                                                  30'd    2895    : data = 32'h    41A5DA13    ;    //    srai x20 x11 26      ====        srai s4, a1, 26
                                                  30'd    2896    : data = 32'h    014D2B33    ;    //    slt x22 x26 x20      ====        slt s6, s10, s4
                                                  30'd    2897    : data = 32'h    01350733    ;    //    add x14 x10 x19      ====        add a4, a0, s3
                                                  30'd    2898    : data = 32'h    09A33613    ;    //    sltiu x12 x6 154      ====        sltiu a2, t1, 154
                                                  30'd    2899    : data = 32'h    3561E4B7    ;    //    lui x9 218654      ====        lui s1, 218654
                                                  30'd    2900    : data = 32'h    43BD0913    ;    //    addi x18 x26 1083      ====        addi s2, s10, 1083
                                                  30'd    2901    : data = 32'h    01BD1493    ;    //    slli x9 x26 27      ====        slli s1, s10, 27
                                                  30'd    2902    : data = 32'h    D51B0713    ;    //    addi x14 x22 -687      ====        addi a4, s6, -687
                                                  30'd    2903    : data = 32'h    F87F4493    ;    //    xori x9 x30 -121      ====        xori s1, t5, -121
                                                  30'd    2904    : data = 32'h    41A80733    ;    //    sub x14 x16 x26      ====        sub a4, a6, s10
                                                  30'd    2905    : data = 32'h    418354B3    ;    //    sra x9 x6 x24      ====        sra s1, t1, s8
                                                  30'd    2906    : data = 32'h    A07A0817    ;    //    auipc x16 657312      ====        auipc a6, 657312
                                                  30'd    2907    : data = 32'h    FECD0897    ;    //    auipc x17 1043664      ====        auipc a7, 1043664
                                                  30'd    2908    : data = 32'h    0160FCB3    ;    //    and x25 x1 x22      ====        and s9, ra, s6
                                                  30'd    2909    : data = 32'h    00E20133    ;    //    add x2 x4 x14      ====        add sp, tp, a4
                                                  30'd    2910    : data = 32'h    8EA16713    ;    //    ori x14 x2 -1814      ====        ori a4, sp, -1814
                                                  30'd    2911    : data = 32'h    001EAA33    ;    //    slt x20 x29 x1      ====        slt s4, t4, ra
                                                  30'd    2912    : data = 32'h    014F55B3    ;    //    srl x11 x30 x20      ====        srl a1, t5, s4
                                                  30'd    2913    : data = 32'h    5FE10817    ;    //    auipc x16 392720      ====        auipc a6, 392720
                                                  30'd    2914    : data = 32'h    01BC8433    ;    //    add x8 x25 x27      ====        add s0, s9, s11
                                                  30'd    2915    : data = 32'h    708E6993    ;    //    ori x19 x28 1800      ====        ori s3, t3, 1800
                                                  30'd    2916    : data = 32'h    0144EA33    ;    //    or x20 x9 x20      ====        or s4, s1, s4
                                                  30'd    2917    : data = 32'h    003B9CB3    ;    //    sll x25 x23 x3      ====        sll s9, s7, gp
                                                  30'd    2918    : data = 32'h    01555E33    ;    //    srl x28 x10 x21      ====        srl t3, a0, s5
                                                  30'd    2919    : data = 32'h    406B0733    ;    //    sub x14 x22 x6      ====        sub a4, s6, t1
                                                  30'd    2920    : data = 32'h    015C1E13    ;    //    slli x28 x24 21      ====        slli t3, s8, 21
                                                  30'd    2921    : data = 32'h    5D86D817    ;    //    auipc x16 383085      ====        auipc a6, 383085
                                                  30'd    2922    : data = 32'h    0069EB33    ;    //    or x22 x19 x6      ====        or s6, s3, t1
                                                  30'd    2923    : data = 32'h    00722733    ;    //    slt x14 x4 x7      ====        slt a4, tp, t2
                                                  30'd    2924    : data = 32'h    FF9E5B17    ;    //    auipc x22 1047013      ====        auipc s6, 1047013
                                                  30'd    2925    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2926    : data = 32'h    013A6633    ;    //    or x12 x20 x19      ====        or a2, s4, s3
                                                  30'd    2927    : data = 32'h    01896D33    ;    //    or x26 x18 x24      ====        or s10, s2, s8
                                                  30'd    2928    : data = 32'h    00D5EB33    ;    //    or x22 x11 x13      ====        or s6, a1, a3
                                                  30'd    2929    : data = 32'h    00C847B3    ;    //    xor x15 x16 x12      ====        xor a5, a6, a2
                                                  30'd    2930    : data = 32'h    006DD193    ;    //    srli x3 x27 6      ====        srli gp, s11, 6
                                                  30'd    2931    : data = 32'h    01D11713    ;    //    slli x14 x2 29      ====        slli a4, sp, 29
                                                  30'd    2932    : data = 32'h    00331C33    ;    //    sll x24 x6 x3      ====        sll s8, t1, gp
                                                  30'd    2933    : data = 32'h    010FDD93    ;    //    srli x27 x31 16      ====        srli s11, t6, 16
                                                  30'd    2934    : data = 32'h    00FEA833    ;    //    slt x16 x29 x15      ====        slt a6, t4, a5
                                                  30'd    2935    : data = 32'h    0007DAB3    ;    //    srl x21 x15 x0      ====        srl s5, a5, zero
                                                  30'd    2936    : data = 32'h    B89E0993    ;    //    addi x19 x28 -1143      ====        addi s3, t3, -1143
                                                  30'd    2937    : data = 32'h    748BFA13    ;    //    andi x20 x23 1864      ====        andi s4, s7, 1864
                                                  30'd    2938    : data = 32'h    41A4D333    ;    //    sra x6 x9 x26      ====        sra t1, s1, s10
                                                  30'd    2939    : data = 32'h    408A80B3    ;    //    sub x1 x21 x8      ====        sub ra, s5, s0
                                                  30'd    2940    : data = 32'h    4DA3F393    ;    //    andi x7 x7 1242      ====        andi t2, t2, 1242
                                                  30'd    2941    : data = 32'h    4186DDB3    ;    //    sra x27 x13 x24      ====        sra s11, a3, s8
                                                  30'd    2942    : data = 32'h    F16CC937    ;    //    lui x18 988876      ====        lui s2, 988876
                                                  30'd    2943    : data = 32'h    007543B3    ;    //    xor x7 x10 x7      ====        xor t2, a0, t2
                                                  30'd    2944    : data = 32'h    CE7EC7B7    ;    //    lui x15 845804      ====        lui a5, 845804
                                                  30'd    2945    : data = 32'h    64D607B7    ;    //    lui x15 413024      ====        lui a5, 413024
                                                  30'd    2946    : data = 32'h    A665CC97    ;    //    auipc x25 681564      ====        auipc s9, 681564
                                                  30'd    2947    : data = 32'h    0172B633    ;    //    sltu x12 x5 x23      ====        sltu a2, t0, s7
                                                  30'd    2948    : data = 32'h    016152B3    ;    //    srl x5 x2 x22      ====        srl t0, sp, s6
                                                  30'd    2949    : data = 32'h    40AA55B3    ;    //    sra x11 x20 x10      ====        sra a1, s4, a0
                                                  30'd    2950    : data = 32'h    B8D96093    ;    //    ori x1 x18 -1139      ====        ori ra, s2, -1139
                                                  30'd    2951    : data = 32'h    4F932417    ;    //    auipc x8 325938      ====        auipc s0, 325938
                                                  30'd    2952    : data = 32'h    4659D937    ;    //    lui x18 288157      ====        lui s2, 288157
                                                  30'd    2953    : data = 32'h    1BE7AC13    ;    //    slti x24 x15 446      ====        slti s8, a5, 446
                                                  30'd    2954    : data = 32'h    403A5F93    ;    //    srai x31 x20 3      ====        srai t6, s4, 3
                                                  30'd    2955    : data = 32'h    01F17B33    ;    //    and x22 x2 x31      ====        and s6, sp, t6
                                                  30'd    2956    : data = 32'h    40B58EB3    ;    //    sub x29 x11 x11      ====        sub t4, a1, a1
                                                  30'd    2957    : data = 32'h    01F20133    ;    //    add x2 x4 x31      ====        add sp, tp, t6
                                                  30'd    2958    : data = 32'h    401A01B3    ;    //    sub x3 x20 x1      ====        sub gp, s4, ra
                                                  30'd    2959    : data = 32'h    FD8E9397    ;    //    auipc x7 1038569      ====        auipc t2, 1038569
                                                  30'd    2960    : data = 32'h    014EA1B3    ;    //    slt x3 x29 x20      ====        slt gp, t4, s4
                                                  30'd    2961    : data = 32'h    00849CB3    ;    //    sll x25 x9 x8      ====        sll s9, s1, s0
                                                  30'd    2962    : data = 32'h    00435613    ;    //    srli x12 x6 4      ====        srli a2, t1, 4
                                                  30'd    2963    : data = 32'h    002BD2B3    ;    //    srl x5 x23 x2      ====        srl t0, s7, sp
                                                  30'd    2964    : data = 32'h    0106D0B3    ;    //    srl x1 x13 x16      ====        srl ra, a3, a6
                                                  30'd    2965    : data = 32'h    636E0097    ;    //    auipc x1 407264      ====        auipc ra, 407264
                                                  30'd    2966    : data = 32'h    0052BEB3    ;    //    sltu x29 x5 x5      ====        sltu t4, t0, t0
                                                  30'd    2967    : data = 32'h    410687B3    ;    //    sub x15 x13 x16      ====        sub a5, a3, a6
                                                  30'd    2968    : data = 32'h    403554B3    ;    //    sra x9 x10 x3      ====        sra s1, a0, gp
                                                  30'd    2969    : data = 32'h    3E887AB7    ;    //    lui x21 256135      ====        lui s5, 256135
                                                  30'd    2970    : data = 32'h    0138AEB3    ;    //    slt x29 x17 x19      ====        slt t4, a7, s3
                                                  30'd    2971    : data = 32'h    3A0D0393    ;    //    addi x7 x26 928      ====        addi t2, s10, 928
                                                  30'd    2972    : data = 32'h    01F689B3    ;    //    add x19 x13 x31      ====        add s3, a3, t6
                                                  30'd    2973    : data = 32'h    4193D633    ;    //    sra x12 x7 x25      ====        sra a2, t2, s9
                                                  30'd    2974    : data = 32'h    6DC5AD13    ;    //    slti x26 x11 1756      ====        slti s10, a1, 1756
                                                  30'd    2975    : data = 32'h    01D3D713    ;    //    srli x14 x7 29      ====        srli a4, t2, 29
                                                  30'd    2976    : data = 32'h    016E39B3    ;    //    sltu x19 x28 x22      ====        sltu s3, t3, s6
                                                  30'd    2977    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    2978    : data = 32'h    41AF02B3    ;    //    sub x5 x30 x26      ====        sub t0, t5, s10
                                                  30'd    2979    : data = 32'h    41F5D2B3    ;    //    sra x5 x11 x31      ====        sra t0, a1, t6
                                                  30'd    2980    : data = 32'h    4124DD93    ;    //    srai x27 x9 18      ====        srai s11, s1, 18
                                                  30'd    2981    : data = 32'h    00939613    ;    //    slli x12 x7 9      ====        slli a2, t2, 9
                                                  30'd    2982    : data = 32'h    01FD3C33    ;    //    sltu x24 x26 x31      ====        sltu s8, s10, t6
                                                  30'd    2983    : data = 32'h    009BADB3    ;    //    slt x27 x23 x9      ====        slt s11, s7, s1
                                                  30'd    2984    : data = 32'h    B705C097    ;    //    auipc x1 749660      ====        auipc ra, 749660
                                                  30'd    2985    : data = 32'h    01CDD133    ;    //    srl x2 x27 x28      ====        srl sp, s11, t3
                                                  30'd    2986    : data = 32'h    019C3833    ;    //    sltu x16 x24 x25      ====        sltu a6, s8, s9
                                                  30'd    2987    : data = 32'h    1A852393    ;    //    slti x7 x10 424      ====        slti t2, a0, 424
                                                  30'd    2988    : data = 32'h    40220933    ;    //    sub x18 x4 x2      ====        sub s2, tp, sp
                                                  30'd    2989    : data = 32'h    DC29B993    ;    //    sltiu x19 x19 -574      ====        sltiu s3, s3, -574
                                                  30'd    2990    : data = 32'h    010261B3    ;    //    or x3 x4 x16      ====        or gp, tp, a6
                                                  30'd    2991    : data = 32'h    018AC633    ;    //    xor x12 x21 x24      ====        xor a2, s5, s8
                                                  30'd    2992    : data = 32'h    017527B3    ;    //    slt x15 x10 x23      ====        slt a5, a0, s7
                                                  30'd    2993    : data = 32'h    401E5D13    ;    //    srai x26 x28 1      ====        srai s10, t3, 1
                                                  30'd    2994    : data = 32'h    B8C86D93    ;    //    ori x27 x16 -1140      ====        ori s11, a6, -1140
                                                  30'd    2995    : data = 32'h    8B78A437    ;    //    lui x8 571274      ====        lui s0, 571274
                                                  30'd    2996    : data = 32'h    404AD833    ;    //    sra x16 x21 x4      ====        sra a6, s5, tp
                                                  30'd    2997    : data = 32'h    00510733    ;    //    add x14 x2 x5      ====        add a4, sp, t0
                                                  30'd    2998    : data = 32'h    006F5913    ;    //    srli x18 x30 6      ====        srli s2, t5, 6
                                                  30'd    2999    : data = 32'h    40945AB3    ;    //    sra x21 x8 x9      ====        sra s5, s0, s1
                                                  30'd    3000    : data = 32'h    331AF4B7    ;    //    lui x9 209327      ====        lui s1, 209327
                                                  30'd    3001    : data = 32'h    01A141B3    ;    //    xor x3 x2 x26      ====        xor gp, sp, s10
                                                  30'd    3002    : data = 32'h    41AD5FB3    ;    //    sra x31 x26 x26      ====        sra t6, s10, s10
                                                  30'd    3003    : data = 32'h    6E15E313    ;    //    ori x6 x11 1761      ====        ori t1, a1, 1761
                                                  30'd    3004    : data = 32'h    005F2B33    ;    //    slt x22 x30 x5      ====        slt s6, t5, t0
                                                  30'd    3005    : data = 32'h    01DD34B3    ;    //    sltu x9 x26 x29      ====        sltu s1, s10, t4
                                                  30'd    3006    : data = 32'h    001F6A33    ;    //    or x20 x30 x1      ====        or s4, t5, ra
                                                  30'd    3007    : data = 32'h    01501B33    ;    //    sll x22 x0 x21      ====        sll s6, zero, s5
                                                  30'd    3008    : data = 32'h    019C35B3    ;    //    sltu x11 x24 x25      ====        sltu a1, s8, s9
                                                  30'd    3009    : data = 32'h    01C8A7B3    ;    //    slt x15 x17 x28      ====        slt a5, a7, t3
                                                  30'd    3010    : data = 32'h    407488B3    ;    //    sub x17 x9 x7      ====        sub a7, s1, t2
                                                  30'd    3011    : data = 32'h    42D8A937    ;    //    lui x18 273802      ====        lui s2, 273802
                                                  30'd    3012    : data = 32'h    40555D13    ;    //    srai x26 x10 5      ====        srai s10, a0, 5
                                                  30'd    3013    : data = 32'h    DFE03893    ;    //    sltiu x17 x0 -514      ====        sltiu a7, zero, -514
                                                  30'd    3014    : data = 32'h    00808E33    ;    //    add x28 x1 x8      ====        add t3, ra, s0
                                                  30'd    3015    : data = 32'h    0175C1B3    ;    //    xor x3 x11 x23      ====        xor gp, a1, s7
                                                  30'd    3016    : data = 32'h    005F2E33    ;    //    slt x28 x30 x5      ====        slt t3, t5, t0
                                                  30'd    3017    : data = 32'h    39F1A593    ;    //    slti x11 x3 927      ====        slti a1, gp, 927
                                                  30'd    3018    : data = 32'h    010A1633    ;    //    sll x12 x20 x16      ====        sll a2, s4, a6
                                                  30'd    3019    : data = 32'h    D9CE6917    ;    //    auipc x18 892134      ====        auipc s2, 892134
                                                  30'd    3020    : data = 32'h    4171DCB3    ;    //    sra x25 x3 x23      ====        sra s9, gp, s7
                                                  30'd    3021    : data = 32'h    055A5397    ;    //    auipc x7 21925      ====        auipc t2, 21925
                                                  30'd    3022    : data = 32'h    0178E9B3    ;    //    or x19 x17 x23      ====        or s3, a7, s7
                                                  30'd    3023    : data = 32'h    0049F833    ;    //    and x16 x19 x4      ====        and a6, s3, tp
                                                  30'd    3024    : data = 32'h    0086DC33    ;    //    srl x24 x13 x8      ====        srl s8, a3, s0
                                                  30'd    3025    : data = 32'h    05ECE613    ;    //    ori x12 x25 94      ====        ori a2, s9, 94
                                                  30'd    3026    : data = 32'h    6673C793    ;    //    xori x15 x7 1639      ====        xori a5, t2, 1639
                                                  30'd    3027    : data = 32'h    0101DE13    ;    //    srli x28 x3 16      ====        srli t3, gp, 16
                                                  30'd    3028    : data = 32'h    40B553B3    ;    //    sra x7 x10 x11      ====        sra t2, a0, a1
                                                  30'd    3029    : data = 32'h    00FC9A13    ;    //    slli x20 x25 15      ====        slli s4, s9, 15
                                                  30'd    3030    : data = 32'h    269673B7    ;    //    lui x7 158055      ====        lui t2, 158055
                                                  30'd    3031    : data = 32'h    015D9493    ;    //    slli x9 x27 21      ====        slli s1, s11, 21
                                                  30'd    3032    : data = 32'h    716BA417    ;    //    auipc x8 464570      ====        auipc s0, 464570
                                                  30'd    3033    : data = 32'h    AFD57713    ;    //    andi x14 x10 -1283      ====        andi a4, a0, -1283
                                                  30'd    3034    : data = 32'h    00974A13    ;    //    xori x20 x14 9      ====        xori s4, a4, 9
                                                  30'd    3035    : data = 32'h    BD5A6B13    ;    //    ori x22 x20 -1067      ====        ori s6, s4, -1067
                                                  30'd    3036    : data = 32'h    010DF9B3    ;    //    and x19 x27 x16      ====        and s3, s11, a6
                                                  30'd    3037    : data = 32'h    6D7AB9B7    ;    //    lui x19 448427      ====        lui s3, 448427
                                                  30'd    3038    : data = 32'h    40C280B3    ;    //    sub x1 x5 x12      ====        sub ra, t0, a2
                                                  30'd    3039    : data = 32'h    00985FB3    ;    //    srl x31 x16 x9      ====        srl t6, a6, s1
                                                  30'd    3040    : data = 32'h    01745913    ;    //    srli x18 x8 23      ====        srli s2, s0, 23
                                                  30'd    3041    : data = 32'h    00E91BB3    ;    //    sll x23 x18 x14      ====        sll s7, s2, a4
                                                  30'd    3042    : data = 32'h    019625B3    ;    //    slt x11 x12 x25      ====        slt a1, a2, s9
                                                  30'd    3043    : data = 32'h    A0B3A5B7    ;    //    lui x11 658234      ====        lui a1, 658234
                                                  30'd    3044    : data = 32'h    0092B733    ;    //    sltu x14 x5 x9      ====        sltu a4, t0, s1
                                                  30'd    3045    : data = 32'h    41D8D593    ;    //    srai x11 x17 29      ====        srai a1, a7, 29
                                                  30'd    3046    : data = 32'h    000189B3    ;    //    add x19 x3 x0      ====        add s3, gp, zero
                                                  30'd    3047    : data = 32'h    01774333    ;    //    xor x6 x14 x23      ====        xor t1, a4, s7
                                                  30'd    3048    : data = 32'h    06680C93    ;    //    addi x25 x16 102      ====        addi s9, a6, 102
                                                  30'd    3049    : data = 32'h    E9717597    ;    //    auipc x11 956183      ====        auipc a1, 956183
                                                  30'd    3050    : data = 32'h    01A1D933    ;    //    srl x18 x3 x26      ====        srl s2, gp, s10
                                                  30'd    3051    : data = 32'h    64F28293    ;    //    addi x5 x5 1615      ====        addi t0, t0, 1615
                                                  30'd    3052    : data = 32'h    EE3C4693    ;    //    xori x13 x24 -285      ====        xori a3, s8, -285
                                                  30'd    3053    : data = 32'h    E2286A13    ;    //    ori x20 x16 -478      ====        ori s4, a6, -478
                                                  30'd    3054    : data = 32'h    5618F713    ;    //    andi x14 x17 1377      ====        andi a4, a7, 1377
                                                  30'd    3055    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3056    : data = 32'h    5A878337    ;    //    lui x6 370808      ====        lui t1, 370808
                                                  30'd    3057    : data = 32'h    4F1FD297    ;    //    auipc x5 324093      ====        auipc t0, 324093
                                                  30'd    3058    : data = 32'h    006078B3    ;    //    and x17 x0 x6      ====        and a7, zero, t1
                                                  30'd    3059    : data = 32'h    5F546E13    ;    //    ori x28 x8 1525      ====        ori t3, s0, 1525
                                                  30'd    3060    : data = 32'h    49A9D797    ;    //    auipc x15 301725      ====        auipc a5, 301725
                                                  30'd    3061    : data = 32'h    DE53FB13    ;    //    andi x22 x7 -539      ====        andi s6, t2, -539
                                                  30'd    3062    : data = 32'h    4103D793    ;    //    srai x15 x7 16      ====        srai a5, t2, 16
                                                  30'd    3063    : data = 32'h    01F87D33    ;    //    and x26 x16 x31      ====        and s10, a6, t6
                                                  30'd    3064    : data = 32'h    0029C333    ;    //    xor x6 x19 x2      ====        xor t1, s3, sp
                                                  30'd    3065    : data = 32'h    003BDE93    ;    //    srli x29 x23 3      ====        srli t4, s7, 3
                                                  30'd    3066    : data = 32'h    003CADB3    ;    //    slt x27 x25 x3      ====        slt s11, s9, gp
                                                  30'd    3067    : data = 32'h    267D6E13    ;    //    ori x28 x26 615      ====        ori t3, s10, 615
                                                  30'd    3068    : data = 32'h    40CAD4B3    ;    //    sra x9 x21 x12      ====        sra s1, s5, a2
                                                  30'd    3069    : data = 32'h    7595CC13    ;    //    xori x24 x11 1881      ====        xori s8, a1, 1881
                                                  30'd    3070    : data = 32'h    76848A93    ;    //    addi x21 x9 1896      ====        addi s5, s1, 1896
                                                  30'd    3071    : data = 32'h    02E15B37    ;    //    lui x22 11797      ====        lui s6, 11797
                                                  30'd    3072    : data = 32'h    B80FB193    ;    //    sltiu x3 x31 -1152      ====        sltiu gp, t6, -1152
                                                  30'd    3073    : data = 32'h    00B00733    ;    //    add x14 x0 x11      ====        add a4, zero, a1
                                                  30'd    3074    : data = 32'h    A7F6C893    ;    //    xori x17 x13 -1409      ====        xori a7, a3, -1409
                                                  30'd    3075    : data = 32'h    01ADE333    ;    //    or x6 x27 x26      ====        or t1, s11, s10
                                                  30'd    3076    : data = 32'h    008DEFB3    ;    //    or x31 x27 x8      ====        or t6, s11, s0
                                                  30'd    3077    : data = 32'h    00EF2AB3    ;    //    slt x21 x30 x14      ====        slt s5, t5, a4
                                                  30'd    3078    : data = 32'h    00E678B3    ;    //    and x17 x12 x14      ====        and a7, a2, a4
                                                  30'd    3079    : data = 32'h    20360613    ;    //    addi x12 x12 515      ====        addi a2, a2, 515
                                                  30'd    3080    : data = 32'h    00BC81B3    ;    //    add x3 x25 x11      ====        add gp, s9, a1
                                                  30'd    3081    : data = 32'h    01F904B3    ;    //    add x9 x18 x31      ====        add s1, s2, t6
                                                  30'd    3082    : data = 32'h    41F95813    ;    //    srai x16 x18 31      ====        srai a6, s2, 31
                                                  30'd    3083    : data = 32'h    0070FE33    ;    //    and x28 x1 x7      ====        and t3, ra, t2
                                                  30'd    3084    : data = 32'h    01BA7B33    ;    //    and x22 x20 x27      ====        and s6, s4, s11
                                                  30'd    3085    : data = 32'h    01DF9A13    ;    //    slli x20 x31 29      ====        slli s4, t6, 29
                                                  30'd    3086    : data = 32'h    41AA06B3    ;    //    sub x13 x20 x26      ====        sub a3, s4, s10
                                                  30'd    3087    : data = 32'h    0290A413    ;    //    slti x8 x1 41      ====        slti s0, ra, 41
                                                  30'd    3088    : data = 32'h    A07C7713    ;    //    andi x14 x24 -1529      ====        andi a4, s8, -1529
                                                  30'd    3089    : data = 32'h    90337413    ;    //    andi x8 x6 -1789      ====        andi s0, t1, -1789
                                                  30'd    3090    : data = 32'h    A63EA897    ;    //    auipc x17 680938      ====        auipc a7, 680938
                                                  30'd    3091    : data = 32'h    93B16597    ;    //    auipc x11 604950      ====        auipc a1, 604950
                                                  30'd    3092    : data = 32'h    01B32CB3    ;    //    slt x25 x6 x27      ====        slt s9, t1, s11
                                                  30'd    3093    : data = 32'h    00DF7D33    ;    //    and x26 x30 x13      ====        and s10, t5, a3
                                                  30'd    3094    : data = 32'h    01CBDBB3    ;    //    srl x23 x23 x28      ====        srl s7, s7, t3
                                                  30'd    3095    : data = 32'h    00A61D33    ;    //    sll x26 x12 x10      ====        sll s10, a2, a0
                                                  30'd    3096    : data = 32'h    403ED313    ;    //    srai x6 x29 3      ====        srai t1, t4, 3
                                                  30'd    3097    : data = 32'h    0119D193    ;    //    srli x3 x19 17      ====        srli gp, s3, 17
                                                  30'd    3098    : data = 32'h    01D4AC33    ;    //    slt x24 x9 x29      ====        slt s8, s1, t4
                                                  30'd    3099    : data = 32'h    342CEE13    ;    //    ori x28 x25 834      ====        ori t3, s9, 834
                                                  30'd    3100    : data = 32'h    A416A617    ;    //    auipc x12 672106      ====        auipc a2, 672106
                                                  30'd    3101    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3102    : data = 32'h    D88F6893    ;    //    ori x17 x30 -632      ====        ori a7, t5, -632
                                                  30'd    3103    : data = 32'h    01617733    ;    //    and x14 x2 x22      ====        and a4, sp, s6
                                                  30'd    3104    : data = 32'h    013AD733    ;    //    srl x14 x21 x19      ====        srl a4, s5, s3
                                                  30'd    3105    : data = 32'h    00AC6333    ;    //    or x6 x24 x10      ====        or t1, s8, a0
                                                  30'd    3106    : data = 32'h    01E2D0B3    ;    //    srl x1 x5 x30      ====        srl ra, t0, t5
                                                  30'd    3107    : data = 32'h    AA470493    ;    //    addi x9 x14 -1372      ====        addi s1, a4, -1372
                                                  30'd    3108    : data = 32'h    01B5CDB3    ;    //    xor x27 x11 x27      ====        xor s11, a1, s11
                                                  30'd    3109    : data = 32'h    B0D16713    ;    //    ori x14 x2 -1267      ====        ori a4, sp, -1267
                                                  30'd    3110    : data = 32'h    004B46B3    ;    //    xor x13 x22 x4      ====        xor a3, s6, tp
                                                  30'd    3111    : data = 32'h    DA6F3293    ;    //    sltiu x5 x30 -602      ====        sltiu t0, t5, -602
                                                  30'd    3112    : data = 32'h    78090113    ;    //    addi x2 x18 1920      ====        addi sp, s2, 1920
                                                  30'd    3113    : data = 32'h    00A3D793    ;    //    srli x15 x7 10      ====        srli a5, t2, 10
                                                  30'd    3114    : data = 32'h    34196C13    ;    //    ori x24 x18 833      ====        ori s8, s2, 833
                                                  30'd    3115    : data = 32'h    39D59137    ;    //    lui x2 236889      ====        lui sp, 236889
                                                  30'd    3116    : data = 32'h    002FDF93    ;    //    srli x31 x31 2      ====        srli t6, t6, 2
                                                  30'd    3117    : data = 32'h    A0514AB7    ;    //    lui x21 656660      ====        lui s5, 656660
                                                  30'd    3118    : data = 32'h    00BEB633    ;    //    sltu x12 x29 x11      ====        sltu a2, t4, a1
                                                  30'd    3119    : data = 32'h    0022F3B3    ;    //    and x7 x5 x2      ====        and t2, t0, sp
                                                  30'd    3120    : data = 32'h    7EE7FA13    ;    //    andi x20 x15 2030      ====        andi s4, a5, 2030
                                                  30'd    3121    : data = 32'h    DFFB4E93    ;    //    xori x29 x22 -513      ====        xori t4, s6, -513
                                                  30'd    3122    : data = 32'h    A6DC8F93    ;    //    addi x31 x25 -1427      ====        addi t6, s9, -1427
                                                  30'd    3123    : data = 32'h    3C4F3693    ;    //    sltiu x13 x30 964      ====        sltiu a3, t5, 964
                                                  30'd    3124    : data = 32'h    013946B3    ;    //    xor x13 x18 x19      ====        xor a3, s2, s3
                                                  30'd    3125    : data = 32'h    012A60B3    ;    //    or x1 x20 x18      ====        or ra, s4, s2
                                                  30'd    3126    : data = 32'h    008B42B3    ;    //    xor x5 x22 x8      ====        xor t0, s6, s0
                                                  30'd    3127    : data = 32'h    016B12B3    ;    //    sll x5 x22 x22      ====        sll t0, s6, s6
                                                  30'd    3128    : data = 32'h    828D3F93    ;    //    sltiu x31 x26 -2008      ====        sltiu t6, s10, -2008
                                                  30'd    3129    : data = 32'h    5A272813    ;    //    slti x16 x14 1442      ====        slti a6, a4, 1442
                                                  30'd    3130    : data = 32'h    2594A493    ;    //    slti x9 x9 601      ====        slti s1, s1, 601
                                                  30'd    3131    : data = 32'h    01810D33    ;    //    add x26 x2 x24      ====        add s10, sp, s8
                                                  30'd    3132    : data = 32'h    1FAFB293    ;    //    sltiu x5 x31 506      ====        sltiu t0, t6, 506
                                                  30'd    3133    : data = 32'h    445E0293    ;    //    addi x5 x28 1093      ====        addi t0, t3, 1093
                                                  30'd    3134    : data = 32'h    00DA19B3    ;    //    sll x19 x20 x13      ====        sll s3, s4, a3
                                                  30'd    3135    : data = 32'h    00792733    ;    //    slt x14 x18 x7      ====        slt a4, s2, t2
                                                  30'd    3136    : data = 32'h    4FF7F613    ;    //    andi x12 x15 1279      ====        andi a2, a5, 1279
                                                  30'd    3137    : data = 32'h    0003ED33    ;    //    or x26 x7 x0      ====        or s10, t2, zero
                                                  30'd    3138    : data = 32'h    37522D13    ;    //    slti x26 x4 885      ====        slti s10, tp, 885
                                                  30'd    3139    : data = 32'h    92C84BB7    ;    //    lui x23 601220      ====        lui s7, 601220
                                                  30'd    3140    : data = 32'h    EC772717    ;    //    auipc x14 968562      ====        auipc a4, 968562
                                                  30'd    3141    : data = 32'h    0112D733    ;    //    srl x14 x5 x17      ====        srl a4, t0, a7
                                                  30'd    3142    : data = 32'h    01F4EA33    ;    //    or x20 x9 x31      ====        or s4, s1, t6
                                                  30'd    3143    : data = 32'h    00B67D33    ;    //    and x26 x12 x11      ====        and s10, a2, a1
                                                  30'd    3144    : data = 32'h    0027B9B3    ;    //    sltu x19 x15 x2      ====        sltu s3, a5, sp
                                                  30'd    3145    : data = 32'h    39806597    ;    //    auipc x11 235526      ====        auipc a1, 235526
                                                  30'd    3146    : data = 32'h    01101893    ;    //    slli x17 x0 17      ====        slli a7, zero, 17
                                                  30'd    3147    : data = 32'h    4C521EB7    ;    //    lui x29 312609      ====        lui t4, 312609
                                                  30'd    3148    : data = 32'h    4A85DB37    ;    //    lui x22 305245      ====        lui s6, 305245
                                                  30'd    3149    : data = 32'h    10AD4813    ;    //    xori x16 x26 266      ====        xori a6, s10, 266
                                                  30'd    3150    : data = 32'h    09B22993    ;    //    slti x19 x4 155      ====        slti s3, tp, 155
                                                  30'd    3151    : data = 32'h    002B8733    ;    //    add x14 x23 x2      ====        add a4, s7, sp
                                                  30'd    3152    : data = 32'h    4BC6A313    ;    //    slti x6 x13 1212      ====        slti t1, a3, 1212
                                                  30'd    3153    : data = 32'h    7C712193    ;    //    slti x3 x2 1991      ====        slti gp, sp, 1991
                                                  30'd    3154    : data = 32'h    001ED3B3    ;    //    srl x7 x29 x1      ====        srl t2, t4, ra
                                                  30'd    3155    : data = 32'h    40085FB3    ;    //    sra x31 x16 x0      ====        sra t6, a6, zero
                                                  30'd    3156    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3157    : data = 32'h    01752D33    ;    //    slt x26 x10 x23      ====        slt s10, a0, s7
                                                  30'd    3158    : data = 32'h    004B5493    ;    //    srli x9 x22 4      ====        srli s1, s6, 4
                                                  30'd    3159    : data = 32'h    40780E33    ;    //    sub x28 x16 x7      ====        sub t3, a6, t2
                                                  30'd    3160    : data = 32'h    5D84F393    ;    //    andi x7 x9 1496      ====        andi t2, s1, 1496
                                                  30'd    3161    : data = 32'h    B6D83813    ;    //    sltiu x16 x16 -1171      ====        sltiu a6, a6, -1171
                                                  30'd    3162    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3163    : data = 32'h    0B1BFE13    ;    //    andi x28 x23 177      ====        andi t3, s7, 177
                                                  30'd    3164    : data = 32'h    FEF78A37    ;    //    lui x20 1044344      ====        lui s4, 1044344
                                                  30'd    3165    : data = 32'h    003FCA33    ;    //    xor x20 x31 x3      ====        xor s4, t6, gp
                                                  30'd    3166    : data = 32'h    01D42733    ;    //    slt x14 x8 x29      ====        slt a4, s0, t4
                                                  30'd    3167    : data = 32'h    008CDD13    ;    //    srli x26 x25 8      ====        srli s10, s9, 8
                                                  30'd    3168    : data = 32'h    010EA833    ;    //    slt x16 x29 x16      ====        slt a6, t4, a6
                                                  30'd    3169    : data = 32'h    B25EE793    ;    //    ori x15 x29 -1243      ====        ori a5, t4, -1243
                                                  30'd    3170    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3171    : data = 32'h    C0323593    ;    //    sltiu x11 x4 -1021      ====        sltiu a1, tp, -1021
                                                  30'd    3172    : data = 32'h    400307B3    ;    //    sub x15 x6 x0      ====        sub a5, t1, zero
                                                  30'd    3173    : data = 32'h    01C643B3    ;    //    xor x7 x12 x28      ====        xor t2, a2, t3
                                                  30'd    3174    : data = 32'h    01B67633    ;    //    and x12 x12 x27      ====        and a2, a2, s11
                                                  30'd    3175    : data = 32'h    11BA19B7    ;    //    lui x19 72609      ====        lui s3, 72609
                                                  30'd    3176    : data = 32'h    D7480813    ;    //    addi x16 x16 -652      ====        addi a6, a6, -652
                                                  30'd    3177    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3178    : data = 32'h    01531033    ;    //    sll x0 x6 x21      ====        sll zero, t1, s5
                                                  30'd    3179    : data = 32'h    00AAD093    ;    //    srli x1 x21 10      ====        srli ra, s5, 10
                                                  30'd    3180    : data = 32'h    4198D593    ;    //    srai x11 x17 25      ====        srai a1, a7, 25
                                                  30'd    3181    : data = 32'h    015A0733    ;    //    add x14 x20 x21      ====        add a4, s4, s5
                                                  30'd    3182    : data = 32'h    0174E433    ;    //    or x8 x9 x23      ====        or s0, s1, s7
                                                  30'd    3183    : data = 32'h    7C95BC13    ;    //    sltiu x24 x11 1993      ====        sltiu s8, a1, 1993
                                                  30'd    3184    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3185    : data = 32'h    AC27A093    ;    //    slti x1 x15 -1342      ====        slti ra, a5, -1342
                                                  30'd    3186    : data = 32'h    008E1433    ;    //    sll x8 x28 x8      ====        sll s0, t3, s0
                                                  30'd    3187    : data = 32'h    7539F493    ;    //    andi x9 x19 1875      ====        andi s1, s3, 1875
                                                  30'd    3188    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3189    : data = 32'h    401C8433    ;    //    sub x8 x25 x1      ====        sub s0, s9, ra
                                                  30'd    3190    : data = 32'h    00BB5EB3    ;    //    srl x29 x22 x11      ====        srl t4, s6, a1
                                                  30'd    3191    : data = 32'h    D566DFB7    ;    //    lui x31 874093      ====        lui t6, 874093
                                                  30'd    3192    : data = 32'h    005FEFB3    ;    //    or x31 x31 x5      ====        or t6, t6, t0
                                                  30'd    3193    : data = 32'h    01C1F2B3    ;    //    and x5 x3 x28      ====        and t0, gp, t3
                                                  30'd    3194    : data = 32'h    019307B3    ;    //    add x15 x6 x25      ====        add a5, t1, s9
                                                  30'd    3195    : data = 32'h    00EE4633    ;    //    xor x12 x28 x14      ====        xor a2, t3, a4
                                                  30'd    3196    : data = 32'h    164F3093    ;    //    sltiu x1 x30 356      ====        sltiu ra, t5, 356
                                                  30'd    3197    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3198    : data = 32'h    6BDBE713    ;    //    ori x14 x23 1725      ====        ori a4, s7, 1725
                                                  30'd    3199    : data = 32'h    1389F193    ;    //    andi x3 x19 312      ====        andi gp, s3, 312
                                                  30'd    3200    : data = 32'h    01854E33    ;    //    xor x28 x10 x24      ====        xor t3, a0, s8
                                                  30'd    3201    : data = 32'h    014B8D33    ;    //    add x26 x23 x20      ====        add s10, s7, s4
                                                  30'd    3202    : data = 32'h    B95A0813    ;    //    addi x16 x20 -1131      ====        addi a6, s4, -1131
                                                  30'd    3203    : data = 32'h    00606DB3    ;    //    or x27 x0 x6      ====        or s11, zero, t1
                                                  30'd    3204    : data = 32'h    018C9713    ;    //    slli x14 x25 24      ====        slli a4, s9, 24
                                                  30'd    3205    : data = 32'h    000ADC13    ;    //    srli x24 x21 0      ====        srli s8, s5, 0
                                                  30'd    3206    : data = 32'h    41FA5413    ;    //    srai x8 x20 31      ====        srai s0, s4, 31
                                                  30'd    3207    : data = 32'h    0074D113    ;    //    srli x2 x9 7      ====        srli sp, s1, 7
                                                  30'd    3208    : data = 32'h    61E30113    ;    //    addi x2 x6 1566      ====        addi sp, t1, 1566
                                                  30'd    3209    : data = 32'h    01339F93    ;    //    slli x31 x7 19      ====        slli t6, t2, 19
                                                  30'd    3210    : data = 32'h    C4F67713    ;    //    andi x14 x12 -945      ====        andi a4, a2, -945
                                                  30'd    3211    : data = 32'h    FD067493    ;    //    andi x9 x12 -48      ====        andi s1, a2, -48
                                                  30'd    3212    : data = 32'h    014376B3    ;    //    and x13 x6 x20      ====        and a3, t1, s4
                                                  30'd    3213    : data = 32'h    01D370B3    ;    //    and x1 x6 x29      ====        and ra, t1, t4
                                                  30'd    3214    : data = 32'h    0003BFB3    ;    //    sltu x31 x7 x0      ====        sltu t6, t2, zero
                                                  30'd    3215    : data = 32'h    C0D58013    ;    //    addi x0 x11 -1011      ====        addi zero, a1, -1011
                                                  30'd    3216    : data = 32'h    011316B3    ;    //    sll x13 x6 x17      ====        sll a3, t1, a7
                                                  30'd    3217    : data = 32'h    C14DC813    ;    //    xori x16 x27 -1004      ====        xori a6, s11, -1004
                                                  30'd    3218    : data = 32'h    6E647B13    ;    //    andi x22 x8 1766      ====        andi s6, s0, 1766
                                                  30'd    3219    : data = 32'h    0046CA33    ;    //    xor x20 x13 x4      ====        xor s4, a3, tp
                                                  30'd    3220    : data = 32'h    01A99793    ;    //    slli x15 x19 26      ====        slli a5, s3, 26
                                                  30'd    3221    : data = 32'h    E9EE6A13    ;    //    ori x20 x28 -354      ====        ori s4, t3, -354
                                                  30'd    3222    : data = 32'h    0038DC33    ;    //    srl x24 x17 x3      ====        srl s8, a7, gp
                                                  30'd    3223    : data = 32'h    504E6A97    ;    //    auipc x21 328934      ====        auipc s5, 328934
                                                  30'd    3224    : data = 32'h    019CF0B3    ;    //    and x1 x25 x25      ====        and ra, s9, s9
                                                  30'd    3225    : data = 32'h    FAF16697    ;    //    auipc x13 1027862      ====        auipc a3, 1027862
                                                  30'd    3226    : data = 32'h    C8EBC593    ;    //    xori x11 x23 -882      ====        xori a1, s7, -882
                                                  30'd    3227    : data = 32'h    01F8E733    ;    //    or x14 x17 x31      ====        or a4, a7, t6
                                                  30'd    3228    : data = 32'h    90814393    ;    //    xori x7 x2 -1784      ====        xori t2, sp, -1784
                                                  30'd    3229    : data = 32'h    402752B3    ;    //    sra x5 x14 x2      ====        sra t0, a4, sp
                                                  30'd    3230    : data = 32'h    78F5A413    ;    //    slti x8 x11 1935      ====        slti s0, a1, 1935
                                                  30'd    3231    : data = 32'h    014AD613    ;    //    srli x12 x21 20      ====        srli a2, s5, 20
                                                  30'd    3232    : data = 32'h    2F976893    ;    //    ori x17 x14 761      ====        ori a7, a4, 761
                                                  30'd    3233    : data = 32'h    01D86DB3    ;    //    or x27 x16 x29      ====        or s11, a6, t4
                                                  30'd    3234    : data = 32'h    00A67BB3    ;    //    and x23 x12 x10      ====        and s7, a2, a0
                                                  30'd    3235    : data = 32'h    003CA2B3    ;    //    slt x5 x25 x3      ====        slt t0, s9, gp
                                                  30'd    3236    : data = 32'h    01B1DBB3    ;    //    srl x23 x3 x27      ====        srl s7, gp, s11
                                                  30'd    3237    : data = 32'h    01DF5033    ;    //    srl x0 x30 x29      ====        srl zero, t5, t4
                                                  30'd    3238    : data = 32'h    1926AC97    ;    //    auipc x25 103018      ====        auipc s9, 103018
                                                  30'd    3239    : data = 32'h    400A86B3    ;    //    sub x13 x21 x0      ====        sub a3, s5, zero
                                                  30'd    3240    : data = 32'h    41DDD013    ;    //    srai x0 x27 29      ====        srai zero, s11, 29
                                                  30'd    3241    : data = 32'h    6136C593    ;    //    xori x11 x13 1555      ====        xori a1, a3, 1555
                                                  30'd    3242    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3243    : data = 32'h    00142AB3    ;    //    slt x21 x8 x1      ====        slt s5, s0, ra
                                                  30'd    3244    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3245    : data = 32'h    41B6DC93    ;    //    srai x25 x13 27      ====        srai s9, a3, 27
                                                  30'd    3246    : data = 32'h    D2053013    ;    //    sltiu x0 x10 -736      ====        sltiu zero, a0, -736
                                                  30'd    3247    : data = 32'h    01E0D813    ;    //    srli x16 x1 30      ====        srli a6, ra, 30
                                                  30'd    3248    : data = 32'h    001E5993    ;    //    srli x19 x28 1      ====        srli s3, t3, 1
                                                  30'd    3249    : data = 32'h    0134F333    ;    //    and x6 x9 x19      ====        and t1, s1, s3
                                                  30'd    3250    : data = 32'h    5F7D0793    ;    //    addi x15 x26 1527      ====        addi a5, s10, 1527
                                                  30'd    3251    : data = 32'h    41495033    ;    //    sra x0 x18 x20      ====        sra zero, s2, s4
                                                  30'd    3252    : data = 32'h    32526693    ;    //    ori x13 x4 805      ====        ori a3, tp, 805
                                                  30'd    3253    : data = 32'h    7368EE17    ;    //    auipc x28 472718      ====        auipc t3, 472718
                                                  30'd    3254    : data = 32'h    01D74DB3    ;    //    xor x27 x14 x29      ====        xor s11, a4, t4
                                                  30'd    3255    : data = 32'h    01EAB333    ;    //    sltu x6 x21 x30      ====        sltu t1, s5, t5
                                                  30'd    3256    : data = 32'h    000F1C93    ;    //    slli x25 x30 0      ====        slli s9, t5, 0
                                                  30'd    3257    : data = 32'h    40668E33    ;    //    sub x28 x13 x6      ====        sub t3, a3, t1
                                                  30'd    3258    : data = 32'h    00644FB3    ;    //    xor x31 x8 x6      ====        xor t6, s0, t1
                                                  30'd    3259    : data = 32'h    64CD2A93    ;    //    slti x21 x26 1612      ====        slti s5, s10, 1612
                                                  30'd    3260    : data = 32'h    407A5393    ;    //    srai x7 x20 7      ====        srai t2, s4, 7
                                                  30'd    3261    : data = 32'h    37EAAB93    ;    //    slti x23 x21 894      ====        slti s7, s5, 894
                                                  30'd    3262    : data = 32'h    00885593    ;    //    srli x11 x16 8      ====        srli a1, a6, 8
                                                  30'd    3263    : data = 32'h    01BAF933    ;    //    and x18 x21 x27      ====        and s2, s5, s11
                                                  30'd    3264    : data = 32'h    407B54B3    ;    //    sra x9 x22 x7      ====        sra s1, s6, t2
                                                  30'd    3265    : data = 32'h    0012AC33    ;    //    slt x24 x5 x1      ====        slt s8, t0, ra
                                                  30'd    3266    : data = 32'h    00BB5093    ;    //    srli x1 x22 11      ====        srli ra, s6, 11
                                                  30'd    3267    : data = 32'h    532BEA93    ;    //    ori x21 x23 1330      ====        ori s5, s7, 1330
                                                  30'd    3268    : data = 32'h    41B688B3    ;    //    sub x17 x13 x27      ====        sub a7, a3, s11
                                                  30'd    3269    : data = 32'h    019CFFB3    ;    //    and x31 x25 x25      ====        and t6, s9, s9
                                                  30'd    3270    : data = 32'h    01620833    ;    //    add x16 x4 x22      ====        add a6, tp, s6
                                                  30'd    3271    : data = 32'h    00C1DD33    ;    //    srl x26 x3 x12      ====        srl s10, gp, a2
                                                  30'd    3272    : data = 32'h    B1708117    ;    //    auipc x2 726792      ====        auipc sp, 726792
                                                  30'd    3273    : data = 32'h    38712F93    ;    //    slti x31 x2 903      ====        slti t6, sp, 903
                                                  30'd    3274    : data = 32'h    E0B34313    ;    //    xori x6 x6 -501      ====        xori t1, t1, -501
                                                  30'd    3275    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3276    : data = 32'h    000C1193    ;    //    slli x3 x24 0      ====        slli gp, s8, 0
                                                  30'd    3277    : data = 32'h    01E3DEB3    ;    //    srl x29 x7 x30      ====        srl t4, t2, t5
                                                  30'd    3278    : data = 32'h    4306EC13    ;    //    ori x24 x13 1072      ====        ori s8, a3, 1072
                                                  30'd    3279    : data = 32'h    00BCD033    ;    //    srl x0 x25 x11      ====        srl zero, s9, a1
                                                  30'd    3280    : data = 32'h    00A1CAB3    ;    //    xor x21 x3 x10      ====        xor s5, gp, a0
                                                  30'd    3281    : data = 32'h    854B3313    ;    //    sltiu x6 x22 -1964      ====        sltiu t1, s6, -1964
                                                  30'd    3282    : data = 32'h    0131B333    ;    //    sltu x6 x3 x19      ====        sltu t1, gp, s3
                                                  30'd    3283    : data = 32'h    40FD8033    ;    //    sub x0 x27 x15      ====        sub zero, s11, a5
                                                  30'd    3284    : data = 32'h    413B5613    ;    //    srai x12 x22 19      ====        srai a2, s6, 19
                                                  30'd    3285    : data = 32'h    00BF48B3    ;    //    xor x17 x30 x11      ====        xor a7, t5, a1
                                                  30'd    3286    : data = 32'h    2B576693    ;    //    ori x13 x14 693      ====        ori a3, a4, 693
                                                  30'd    3287    : data = 32'h    01312033    ;    //    slt x0 x2 x19      ====        slt zero, sp, s3
                                                  30'd    3288    : data = 32'h    017B5D13    ;    //    srli x26 x22 23      ====        srli s10, s6, 23
                                                  30'd    3289    : data = 32'h    F5F9BE17    ;    //    auipc x28 1007515      ====        auipc t3, 1007515
                                                  30'd    3290    : data = 32'h    019ED693    ;    //    srli x13 x29 25      ====        srli a3, t4, 25
                                                  30'd    3291    : data = 32'h    003BF9B3    ;    //    and x19 x23 x3      ====        and s3, s7, gp
                                                  30'd    3292    : data = 32'h    46C53313    ;    //    sltiu x6 x10 1132      ====        sltiu t1, a0, 1132
                                                  30'd    3293    : data = 32'h    402F8D33    ;    //    sub x26 x31 x2      ====        sub s10, t6, sp
                                                  30'd    3294    : data = 32'h    74806D93    ;    //    ori x27 x0 1864      ====        ori s11, zero, 1864
                                                  30'd    3295    : data = 32'h    CCB70E13    ;    //    addi x28 x14 -821      ====        addi t3, a4, -821
                                                  30'd    3296    : data = 32'h    02AA3BB7    ;    //    lui x23 10915      ====        lui s7, 10915
                                                  30'd    3297    : data = 32'h    01DA2733    ;    //    slt x14 x20 x29      ====        slt a4, s4, t4
                                                  30'd    3298    : data = 32'h    00356C33    ;    //    or x24 x10 x3      ====        or s8, a0, gp
                                                  30'd    3299    : data = 32'h    01DB8933    ;    //    add x18 x23 x29      ====        add s2, s7, t4
                                                  30'd    3300    : data = 32'h    66484093    ;    //    xori x1 x16 1636      ====        xori ra, a6, 1636
                                                  30'd    3301    : data = 32'h    78906093    ;    //    ori x1 x0 1929      ====        ori ra, zero, 1929
                                                  30'd    3302    : data = 32'h    00997833    ;    //    and x16 x18 x9      ====        and a6, s2, s1
                                                  30'd    3303    : data = 32'h    00EAC1B3    ;    //    xor x3 x21 x14      ====        xor gp, s5, a4
                                                  30'd    3304    : data = 32'h    007D9933    ;    //    sll x18 x27 x7      ====        sll s2, s11, t2
                                                  30'd    3305    : data = 32'h    CB522013    ;    //    slti x0 x4 -843      ====        slti zero, tp, -843
                                                  30'd    3306    : data = 32'h    003CD113    ;    //    srli x2 x25 3      ====        srli sp, s9, 3
                                                  30'd    3307    : data = 32'h    76803593    ;    //    sltiu x11 x0 1896      ====        sltiu a1, zero, 1896
                                                  30'd    3308    : data = 32'h    006DA333    ;    //    slt x6 x27 x6      ====        slt t1, s11, t1
                                                  30'd    3309    : data = 32'h    DA0DE2B7    ;    //    lui x5 893150      ====        lui t0, 893150
                                                  30'd    3310    : data = 32'h    417C5E93    ;    //    srai x29 x24 23      ====        srai t4, s8, 23
                                                  30'd    3311    : data = 32'h    000111B3    ;    //    sll x3 x2 x0      ====        sll gp, sp, zero
                                                  30'd    3312    : data = 32'h    8B016497    ;    //    auipc x9 569366      ====        auipc s1, 569366
                                                  30'd    3313    : data = 32'h    00502CB3    ;    //    slt x25 x0 x5      ====        slt s9, zero, t0
                                                  30'd    3314    : data = 32'h    40E4DDB3    ;    //    sra x27 x9 x14      ====        sra s11, s1, a4
                                                  30'd    3315    : data = 32'h    00567E33    ;    //    and x28 x12 x5      ====        and t3, a2, t0
                                                  30'd    3316    : data = 32'h    9D244593    ;    //    xori x11 x8 -1582      ====        xori a1, s0, -1582
                                                  30'd    3317    : data = 32'h    6E594C93    ;    //    xori x25 x18 1765      ====        xori s9, s2, 1765
                                                  30'd    3318    : data = 32'h    01331E33    ;    //    sll x28 x6 x19      ====        sll t3, t1, s3
                                                  30'd    3319    : data = 32'h    0C237413    ;    //    andi x8 x6 194      ====        andi s0, t1, 194
                                                  30'd    3320    : data = 32'h    000C1CB3    ;    //    sll x25 x24 x0      ====        sll s9, s8, zero
                                                  30'd    3321    : data = 32'h    00B75433    ;    //    srl x8 x14 x11      ====        srl s0, a4, a1
                                                  30'd    3322    : data = 32'h    1B724613    ;    //    xori x12 x4 439      ====        xori a2, tp, 439
                                                  30'd    3323    : data = 32'h    4022DE13    ;    //    srai x28 x5 2      ====        srai t3, t0, 2
                                                  30'd    3324    : data = 32'h    409DD293    ;    //    srai x5 x27 9      ====        srai t0, s11, 9
                                                  30'd    3325    : data = 32'h    006D2633    ;    //    slt x12 x26 x6      ====        slt a2, s10, t1
                                                  30'd    3326    : data = 32'h    906A6293    ;    //    ori x5 x20 -1786      ====        ori t0, s4, -1786
                                                  30'd    3327    : data = 32'h    405601B3    ;    //    sub x3 x12 x5      ====        sub gp, a2, t0
                                                  30'd    3328    : data = 32'h    41EE57B3    ;    //    sra x15 x28 x30      ====        sra a5, t3, t5
                                                  30'd    3329    : data = 32'h    002F02B3    ;    //    add x5 x30 x2      ====        add t0, t5, sp
                                                  30'd    3330    : data = 32'h    004D0A33    ;    //    add x20 x26 x4      ====        add s4, s10, tp
                                                  30'd    3331    : data = 32'h    007F1A33    ;    //    sll x20 x30 x7      ====        sll s4, t5, t2
                                                  30'd    3332    : data = 32'h    823ED397    ;    //    auipc x7 533485      ====        auipc t2, 533485
                                                  30'd    3333    : data = 32'h    40CDD0B3    ;    //    sra x1 x27 x12      ====        sra ra, s11, a2
                                                  30'd    3334    : data = 32'h    01DB5193    ;    //    srli x3 x22 29      ====        srli gp, s6, 29
                                                  30'd    3335    : data = 32'h    5AEE3A13    ;    //    sltiu x20 x28 1454      ====        sltiu s4, t3, 1454
                                                  30'd    3336    : data = 32'h    4047D833    ;    //    sra x16 x15 x4      ====        sra a6, a5, tp
                                                  30'd    3337    : data = 32'h    542CF313    ;    //    andi x6 x25 1346      ====        andi t1, s9, 1346
                                                  30'd    3338    : data = 32'h    017D1A93    ;    //    slli x21 x26 23      ====        slli s5, s10, 23
                                                  30'd    3339    : data = 32'h    41A151B3    ;    //    sra x3 x2 x26      ====        sra gp, sp, s10
                                                  30'd    3340    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3341    : data = 32'h    41A4DE13    ;    //    srai x28 x9 26      ====        srai t3, s1, 26
                                                  30'd    3342    : data = 32'h    37AE8EB7    ;    //    lui x29 228072      ====        lui t4, 228072
                                                  30'd    3343    : data = 32'h    00195733    ;    //    srl x14 x18 x1      ====        srl a4, s2, ra
                                                  30'd    3344    : data = 32'h    766A0D17    ;    //    auipc x26 485024      ====        auipc s10, 485024
                                                  30'd    3345    : data = 32'h    31667293    ;    //    andi x5 x12 790      ====        andi t0, a2, 790
                                                  30'd    3346    : data = 32'h    40ACDB13    ;    //    srai x22 x25 10      ====        srai s6, s9, 10
                                                  30'd    3347    : data = 32'h    015BBFB3    ;    //    sltu x31 x23 x21      ====        sltu t6, s7, s5
                                                  30'd    3348    : data = 32'h    41E9D7B3    ;    //    sra x15 x19 x30      ====        sra a5, s3, t5
                                                  30'd    3349    : data = 32'h    8A1E2913    ;    //    slti x18 x28 -1887      ====        slti s2, t3, -1887
                                                  30'd    3350    : data = 32'h    013C9913    ;    //    slli x18 x25 19      ====        slli s2, s9, 19
                                                  30'd    3351    : data = 32'h    013C5113    ;    //    srli x2 x24 19      ====        srli sp, s8, 19
                                                  30'd    3352    : data = 32'h    6982B313    ;    //    sltiu x6 x5 1688      ====        sltiu t1, t0, 1688
                                                  30'd    3353    : data = 32'h    D4A74913    ;    //    xori x18 x14 -694      ====        xori s2, a4, -694
                                                  30'd    3354    : data = 32'h    01E6C2B3    ;    //    xor x5 x13 x30      ====        xor t0, a3, t5
                                                  30'd    3355    : data = 32'h    0078D1B3    ;    //    srl x3 x17 x7      ====        srl gp, a7, t2
                                                  30'd    3356    : data = 32'h    03577E93    ;    //    andi x29 x14 53      ====        andi t4, a4, 53
                                                  30'd    3357    : data = 32'h    825BC0B7    ;    //    lui x1 533948      ====        lui ra, 533948
                                                  30'd    3358    : data = 32'h    000C5EB3    ;    //    srl x29 x24 x0      ====        srl t4, s8, zero
                                                  30'd    3359    : data = 32'h    653F6993    ;    //    ori x19 x30 1619      ====        ori s3, t5, 1619
                                                  30'd    3360    : data = 32'h    004948B3    ;    //    xor x17 x18 x4      ====        xor a7, s2, tp
                                                  30'd    3361    : data = 32'h    01F348B3    ;    //    xor x17 x6 x31      ====        xor a7, t1, t6
                                                  30'd    3362    : data = 32'h    18E3AA13    ;    //    slti x20 x7 398      ====        slti s4, t2, 398
                                                  30'd    3363    : data = 32'h    01D1BA33    ;    //    sltu x20 x3 x29      ====        sltu s4, gp, t4
                                                  30'd    3364    : data = 32'h    00D825B3    ;    //    slt x11 x16 x13      ====        slt a1, a6, a3
                                                  30'd    3365    : data = 32'h    B954A1B7    ;    //    lui x3 759114      ====        lui gp, 759114
                                                  30'd    3366    : data = 32'h    5A0FE2B7    ;    //    lui x5 368894      ====        lui t0, 368894
                                                  30'd    3367    : data = 32'h    00CE1933    ;    //    sll x18 x28 x12      ====        sll s2, t3, a2
                                                  30'd    3368    : data = 32'h    016E4A33    ;    //    xor x20 x28 x22      ====        xor s4, t3, s6
                                                  30'd    3369    : data = 32'h    60B4F993    ;    //    andi x19 x9 1547      ====        andi s3, s1, 1547
                                                  30'd    3370    : data = 32'h    0041BDB3    ;    //    sltu x27 x3 x4      ====        sltu s11, gp, tp
                                                  30'd    3371    : data = 32'h    1B787813    ;    //    andi x16 x16 439      ====        andi a6, a6, 439
                                                  30'd    3372    : data = 32'h    011D77B3    ;    //    and x15 x26 x17      ====        and a5, s10, a7
                                                  30'd    3373    : data = 32'h    8D9BF113    ;    //    andi x2 x23 -1831      ====        andi sp, s7, -1831
                                                  30'd    3374    : data = 32'h    0050FA33    ;    //    and x20 x1 x5      ====        and s4, ra, t0
                                                  30'd    3375    : data = 32'h    0008F2B3    ;    //    and x5 x17 x0      ====        and t0, a7, zero
                                                  30'd    3376    : data = 32'h    00B71193    ;    //    slli x3 x14 11      ====        slli gp, a4, 11
                                                  30'd    3377    : data = 32'h    40448833    ;    //    sub x16 x9 x4      ====        sub a6, s1, tp
                                                  30'd    3378    : data = 32'h    3B81E393    ;    //    ori x7 x3 952      ====        ori t2, gp, 952
                                                  30'd    3379    : data = 32'h    00E09113    ;    //    slli x2 x1 14      ====        slli sp, ra, 14
                                                  30'd    3380    : data = 32'h    00FE64B3    ;    //    or x9 x28 x15      ====        or s1, t3, a5
                                                  30'd    3381    : data = 32'h    413858B3    ;    //    sra x17 x16 x19      ====        sra a7, a6, s3
                                                  30'd    3382    : data = 32'h    00FC1933    ;    //    sll x18 x24 x15      ====        sll s2, s8, a5
                                                  30'd    3383    : data = 32'h    CD397E93    ;    //    andi x29 x18 -813      ====        andi t4, s2, -813
                                                  30'd    3384    : data = 32'h    5FC98F93    ;    //    addi x31 x19 1532      ====        addi t6, s3, 1532
                                                  30'd    3385    : data = 32'h    004ADD93    ;    //    srli x27 x21 4      ====        srli s11, s5, 4
                                                  30'd    3386    : data = 32'h    8E18FD13    ;    //    andi x26 x17 -1823      ====        andi s10, a7, -1823
                                                  30'd    3387    : data = 32'h    6D547897    ;    //    auipc x17 447815      ====        auipc a7, 447815
                                                  30'd    3388    : data = 32'h    00A91BB3    ;    //    sll x23 x18 x10      ====        sll s7, s2, a0
                                                  30'd    3389    : data = 32'h    01059E33    ;    //    sll x28 x11 x16      ====        sll t3, a1, a6
                                                  30'd    3390    : data = 32'h    009198B3    ;    //    sll x17 x3 x9      ====        sll a7, gp, s1
                                                  30'd    3391    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3392    : data = 32'h    4145DE33    ;    //    sra x28 x11 x20      ====        sra t3, a1, s4
                                                  30'd    3393    : data = 32'h    011DF333    ;    //    and x6 x27 x17      ====        and t1, s11, a7
                                                  30'd    3394    : data = 32'h    66F32A93    ;    //    slti x21 x6 1647      ====        slti s5, t1, 1647
                                                  30'd    3395    : data = 32'h    97220393    ;    //    addi x7 x4 -1678      ====        addi t2, tp, -1678
                                                  30'd    3396    : data = 32'h    010273B3    ;    //    and x7 x4 x16      ====        and t2, tp, a6
                                                  30'd    3397    : data = 32'h    007710B3    ;    //    sll x1 x14 x7      ====        sll ra, a4, t2
                                                  30'd    3398    : data = 32'h    01DE3A33    ;    //    sltu x20 x28 x29      ====        sltu s4, t3, t4
                                                  30'd    3399    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3400    : data = 32'h    41B7D133    ;    //    sra x2 x15 x27      ====        sra sp, a5, s11
                                                  30'd    3401    : data = 32'h    DE485337    ;    //    lui x6 910469      ====        lui t1, 910469
                                                  30'd    3402    : data = 32'h    408E5A13    ;    //    srai x20 x28 8      ====        srai s4, t3, 8
                                                  30'd    3403    : data = 32'h    000DA433    ;    //    slt x8 x27 x0      ====        slt s0, s11, zero
                                                  30'd    3404    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3405    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3406    : data = 32'h    40485A33    ;    //    sra x20 x16 x4      ====        sra s4, a6, tp
                                                  30'd    3407    : data = 32'h    0DE30413    ;    //    addi x8 x6 222      ====        addi s0, t1, 222
                                                  30'd    3408    : data = 32'h    00D7C133    ;    //    xor x2 x15 x13      ====        xor sp, a5, a3
                                                  30'd    3409    : data = 32'h    01720433    ;    //    add x8 x4 x23      ====        add s0, tp, s7
                                                  30'd    3410    : data = 32'h    DACAB093    ;    //    sltiu x1 x21 -596      ====        sltiu ra, s5, -596
                                                  30'd    3411    : data = 32'h    4A998093    ;    //    addi x1 x19 1193      ====        addi ra, s3, 1193
                                                  30'd    3412    : data = 32'h    00486433    ;    //    or x8 x16 x4      ====        or s0, a6, tp
                                                  30'd    3413    : data = 32'h    008902B3    ;    //    add x5 x18 x8      ====        add t0, s2, s0
                                                  30'd    3414    : data = 32'h    008BA4B3    ;    //    slt x9 x23 x8      ====        slt s1, s7, s0
                                                  30'd    3415    : data = 32'h    008C03B3    ;    //    add x7 x24 x8      ====        add t2, s8, s0
                                                  30'd    3416    : data = 32'h    41935CB3    ;    //    sra x25 x6 x25      ====        sra s9, t1, s9
                                                  30'd    3417    : data = 32'h    41B90633    ;    //    sub x12 x18 x27      ====        sub a2, s2, s11
                                                  30'd    3418    : data = 32'h    00581F93    ;    //    slli x31 x16 5      ====        slli t6, a6, 5
                                                  30'd    3419    : data = 32'h    004F81B3    ;    //    add x3 x31 x4      ====        add gp, t6, tp
                                                  30'd    3420    : data = 32'h    0057DA13    ;    //    srli x20 x15 5      ====        srli s4, a5, 5
                                                  30'd    3421    : data = 32'h    01D60D33    ;    //    add x26 x12 x29      ====        add s10, a2, t4
                                                  30'd    3422    : data = 32'h    3FDA6A37    ;    //    lui x20 261542      ====        lui s4, 261542
                                                  30'd    3423    : data = 32'h    9B0EB893    ;    //    sltiu x17 x29 -1616      ====        sltiu a7, t4, -1616
                                                  30'd    3424    : data = 32'h    406E0833    ;    //    sub x16 x28 x6      ====        sub a6, t3, t1
                                                  30'd    3425    : data = 32'h    FCF7B197    ;    //    auipc x3 1036155      ====        auipc gp, 1036155
                                                  30'd    3426    : data = 32'h    87FB8737    ;    //    lui x14 556984      ====        lui a4, 556984
                                                  30'd    3427    : data = 32'h    0124D893    ;    //    srli x17 x9 18      ====        srli a7, s1, 18
                                                  30'd    3428    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3429    : data = 32'h    CF75B937    ;    //    lui x18 849755      ====        lui s2, 849755
                                                  30'd    3430    : data = 32'h    2C13BE13    ;    //    sltiu x28 x7 705      ====        sltiu t3, t2, 705
                                                  30'd    3431    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3432    : data = 32'h    D12C2D13    ;    //    slti x26 x24 -750      ====        slti s10, s8, -750
                                                  30'd    3433    : data = 32'h    001452B3    ;    //    srl x5 x8 x1      ====        srl t0, s0, ra
                                                  30'd    3434    : data = 32'h    00425633    ;    //    srl x12 x4 x4      ====        srl a2, tp, tp
                                                  30'd    3435    : data = 32'h    003D4BB3    ;    //    xor x23 x26 x3      ====        xor s7, s10, gp
                                                  30'd    3436    : data = 32'h    00745833    ;    //    srl x16 x8 x7      ====        srl a6, s0, t2
                                                  30'd    3437    : data = 32'h    6015C093    ;    //    xori x1 x11 1537      ====        xori ra, a1, 1537
                                                  30'd    3438    : data = 32'h    0133D313    ;    //    srli x6 x7 19      ====        srli t1, t2, 19
                                                  30'd    3439    : data = 32'h    418889B3    ;    //    sub x19 x17 x24      ====        sub s3, a7, s8
                                                  30'd    3440    : data = 32'h    1A9C6B93    ;    //    ori x23 x24 425      ====        ori s7, s8, 425
                                                  30'd    3441    : data = 32'h    79B95797    ;    //    auipc x15 498581      ====        auipc a5, 498581
                                                  30'd    3442    : data = 32'h    006295B3    ;    //    sll x11 x5 x6      ====        sll a1, t0, t1
                                                  30'd    3443    : data = 32'h    A300E313    ;    //    ori x6 x1 -1488      ====        ori t1, ra, -1488
                                                  30'd    3444    : data = 32'h    40B5D133    ;    //    sra x2 x11 x11      ====        sra sp, a1, a1
                                                  30'd    3445    : data = 32'h    00405E93    ;    //    srli x29 x0 4      ====        srli t4, zero, 4
                                                  30'd    3446    : data = 32'h    008B1893    ;    //    slli x17 x22 8      ====        slli a7, s6, 8
                                                  30'd    3447    : data = 32'h    0115A733    ;    //    slt x14 x11 x17      ====        slt a4, a1, a7
                                                  30'd    3448    : data = 32'h    D237E793    ;    //    ori x15 x15 -733      ====        ori a5, a5, -733
                                                  30'd    3449    : data = 32'h    012D78B3    ;    //    and x17 x26 x18      ====        and a7, s10, s2
                                                  30'd    3450    : data = 32'h    407ADEB3    ;    //    sra x29 x21 x7      ====        sra t4, s5, t2
                                                  30'd    3451    : data = 32'h    4133D2B3    ;    //    sra x5 x7 x19      ====        sra t0, t2, s3
                                                  30'd    3452    : data = 32'h    48618D13    ;    //    addi x26 x3 1158      ====        addi s10, gp, 1158
                                                  30'd    3453    : data = 32'h    E9DECD13    ;    //    xori x26 x29 -355      ====        xori s10, t4, -355
                                                  30'd    3454    : data = 32'h    011D5833    ;    //    srl x16 x26 x17      ====        srl a6, s10, a7
                                                  30'd    3455    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3456    : data = 32'h    0626A013    ;    //    slti x0 x13 98      ====        slti zero, a3, 98
                                                  30'd    3457    : data = 32'h    20037693    ;    //    andi x13 x6 512      ====        andi a3, t1, 512
                                                  30'd    3458    : data = 32'h    D861BAB7    ;    //    lui x21 886299      ====        lui s5, 886299
                                                  30'd    3459    : data = 32'h    01CB5393    ;    //    srli x7 x22 28      ====        srli t2, s6, 28
                                                  30'd    3460    : data = 32'h    018723B3    ;    //    slt x7 x14 x24      ====        slt t2, a4, s8
                                                  30'd    3461    : data = 32'h    00EE1893    ;    //    slli x17 x28 14      ====        slli a7, t3, 14
                                                  30'd    3462    : data = 32'h    01E1D113    ;    //    srli x2 x3 30      ====        srli sp, gp, 30
                                                  30'd    3463    : data = 32'h    8C836D37    ;    //    lui x26 575542      ====        lui s10, 575542
                                                  30'd    3464    : data = 32'h    0105DD33    ;    //    srl x26 x11 x16      ====        srl s10, a1, a6
                                                  30'd    3465    : data = 32'h    418CDC33    ;    //    sra x24 x25 x24      ====        sra s8, s9, s8
                                                  30'd    3466    : data = 32'h    DBC0FD13    ;    //    andi x26 x1 -580      ====        andi s10, ra, -580
                                                  30'd    3467    : data = 32'h    007087B3    ;    //    add x15 x1 x7      ====        add a5, ra, t2
                                                  30'd    3468    : data = 32'h    009F9B93    ;    //    slli x23 x31 9      ====        slli s7, t6, 9
                                                  30'd    3469    : data = 32'h    41EF5333    ;    //    sra x6 x30 x30      ====        sra t1, t5, t5
                                                  30'd    3470    : data = 32'h    629BC993    ;    //    xori x19 x23 1577      ====        xori s3, s7, 1577
                                                  30'd    3471    : data = 32'h    17BCCC93    ;    //    xori x25 x25 379      ====        xori s9, s9, 379
                                                  30'd    3472    : data = 32'h    40165313    ;    //    srai x6 x12 1      ====        srai t1, a2, 1
                                                  30'd    3473    : data = 32'h    B41BE113    ;    //    ori x2 x23 -1215      ====        ori sp, s7, -1215
                                                  30'd    3474    : data = 32'h    01B2F8B3    ;    //    and x17 x5 x27      ====        and a7, t0, s11
                                                  30'd    3475    : data = 32'h    01CEC833    ;    //    xor x16 x29 x28      ====        xor a6, t4, t3
                                                  30'd    3476    : data = 32'h    40B28833    ;    //    sub x16 x5 x11      ====        sub a6, t0, a1
                                                  30'd    3477    : data = 32'h    39A86893    ;    //    ori x17 x16 922      ====        ori a7, a6, 922
                                                  30'd    3478    : data = 32'h    F682C293    ;    //    xori x5 x5 -152      ====        xori t0, t0, -152
                                                  30'd    3479    : data = 32'h    F25F9997    ;    //    auipc x19 992761      ====        auipc s3, 992761
                                                  30'd    3480    : data = 32'h    017FD613    ;    //    srli x12 x31 23      ====        srli a2, t6, 23
                                                  30'd    3481    : data = 32'h    01A2DDB3    ;    //    srl x27 x5 x26      ====        srl s11, t0, s10
                                                  30'd    3482    : data = 32'h    404BD433    ;    //    sra x8 x23 x4      ====        sra s0, s7, tp
                                                  30'd    3483    : data = 32'h    22490593    ;    //    addi x11 x18 548      ====        addi a1, s2, 548
                                                  30'd    3484    : data = 32'h    01D5DA93    ;    //    srli x21 x11 29      ====        srli s5, a1, 29
                                                  30'd    3485    : data = 32'h    5C8F8813    ;    //    addi x16 x31 1480      ====        addi a6, t6, 1480
                                                  30'd    3486    : data = 32'h    348E0813    ;    //    addi x16 x28 840      ====        addi a6, t3, 840
                                                  30'd    3487    : data = 32'h    00C751B3    ;    //    srl x3 x14 x12      ====        srl gp, a4, a2
                                                  30'd    3488    : data = 32'h    8B372113    ;    //    slti x2 x14 -1869      ====        slti sp, a4, -1869
                                                  30'd    3489    : data = 32'h    00A9FB33    ;    //    and x22 x19 x10      ====        and s6, s3, a0
                                                  30'd    3490    : data = 32'h    01E11D13    ;    //    slli x26 x2 30      ====        slli s10, sp, 30
                                                  30'd    3491    : data = 32'h    0125ED33    ;    //    or x26 x11 x18      ====        or s10, a1, s2
                                                  30'd    3492    : data = 32'h    00475CB3    ;    //    srl x25 x14 x4      ====        srl s9, a4, tp
                                                  30'd    3493    : data = 32'h    41200AB3    ;    //    sub x21 x0 x18      ====        sub s5, zero, s2
                                                  30'd    3494    : data = 32'h    01CE1DB3    ;    //    sll x27 x28 x28      ====        sll s11, t3, t3
                                                  30'd    3495    : data = 32'h    009C82B3    ;    //    add x5 x25 x9      ====        add t0, s9, s1
                                                  30'd    3496    : data = 32'h    CA0B6017    ;    //    auipc x0 827574      ====        auipc zero, 827574
                                                  30'd    3497    : data = 32'h    A6F8B197    ;    //    auipc x3 683915      ====        auipc gp, 683915
                                                  30'd    3498    : data = 32'h    1C6C8413    ;    //    addi x8 x25 454      ====        addi s0, s9, 454
                                                  30'd    3499    : data = 32'h    D8935137    ;    //    lui x2 887093      ====        lui sp, 887093
                                                  30'd    3500    : data = 32'h    01E0B433    ;    //    sltu x8 x1 x30      ====        sltu s0, ra, t5
                                                  30'd    3501    : data = 32'h    419155B3    ;    //    sra x11 x2 x25      ====        sra a1, sp, s9
                                                  30'd    3502    : data = 32'h    7EBC3A93    ;    //    sltiu x21 x24 2027      ====        sltiu s5, s8, 2027
                                                  30'd    3503    : data = 32'h    3E1953B7    ;    //    lui x7 254357      ====        lui t2, 254357
                                                  30'd    3504    : data = 32'h    00C78DB3    ;    //    add x27 x15 x12      ====        add s11, a5, a2
                                                  30'd    3505    : data = 32'h    2D710A37    ;    //    lui x20 186128      ====        lui s4, 186128
                                                  30'd    3506    : data = 32'h    4180DA33    ;    //    sra x20 x1 x24      ====        sra s4, ra, s8
                                                  30'd    3507    : data = 32'h    E0AAAD13    ;    //    slti x26 x21 -502      ====        slti s10, s5, -502
                                                  30'd    3508    : data = 32'h    CCFD3E13    ;    //    sltiu x28 x26 -817      ====        sltiu t3, s10, -817
                                                  30'd    3509    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3510    : data = 32'h    011126B3    ;    //    slt x13 x2 x17      ====        slt a3, sp, a7
                                                  30'd    3511    : data = 32'h    4051DC33    ;    //    sra x24 x3 x5      ====        sra s8, gp, t0
                                                  30'd    3512    : data = 32'h    3F8D6313    ;    //    ori x6 x26 1016      ====        ori t1, s10, 1016
                                                  30'd    3513    : data = 32'h    00DC9E13    ;    //    slli x28 x25 13      ====        slli t3, s9, 13
                                                  30'd    3514    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3515    : data = 32'h    00B3D7B3    ;    //    srl x15 x7 x11      ====        srl a5, t2, a1
                                                  30'd    3516    : data = 32'h    4AEA6113    ;    //    ori x2 x20 1198      ====        ori sp, s4, 1198
                                                  30'd    3517    : data = 32'h    41C05993    ;    //    srai x19 x0 28      ====        srai s3, zero, 28
                                                  30'd    3518    : data = 32'h    00F11B33    ;    //    sll x22 x2 x15      ====        sll s6, sp, a5
                                                  30'd    3519    : data = 32'h    94832E93    ;    //    slti x29 x6 -1720      ====        slti t4, t1, -1720
                                                  30'd    3520    : data = 32'h    0053D413    ;    //    srli x8 x7 5      ====        srli s0, t2, 5
                                                  30'd    3521    : data = 32'h    010D0733    ;    //    add x14 x26 x16      ====        add a4, s10, a6
                                                  30'd    3522    : data = 32'h    00BF46B3    ;    //    xor x13 x30 x11      ====        xor a3, t5, a1
                                                  30'd    3523    : data = 32'h    016969B3    ;    //    or x19 x18 x22      ====        or s3, s2, s6
                                                  30'd    3524    : data = 32'h    CD254413    ;    //    xori x8 x10 -814      ====        xori s0, a0, -814
                                                  30'd    3525    : data = 32'h    00FEAAB3    ;    //    slt x21 x29 x15      ====        slt s5, t4, a5
                                                  30'd    3526    : data = 32'h    E0AEB013    ;    //    sltiu x0 x29 -502      ====        sltiu zero, t4, -502
                                                  30'd    3527    : data = 32'h    00439A33    ;    //    sll x20 x7 x4      ====        sll s4, t2, tp
                                                  30'd    3528    : data = 32'h    00F97D33    ;    //    and x26 x18 x15      ====        and s10, s2, a5
                                                  30'd    3529    : data = 32'h    01284333    ;    //    xor x6 x16 x18      ====        xor t1, a6, s2
                                                  30'd    3530    : data = 32'h    419DD593    ;    //    srai x11 x27 25      ====        srai a1, s11, 25
                                                  30'd    3531    : data = 32'h    C8F50A13    ;    //    addi x20 x10 -881      ====        addi s4, a0, -881
                                                  30'd    3532    : data = 32'h    00437FB3    ;    //    and x31 x6 x4      ====        and t6, t1, tp
                                                  30'd    3533    : data = 32'h    01EF78B3    ;    //    and x17 x30 x30      ====        and a7, t5, t5
                                                  30'd    3534    : data = 32'h    01B43EB3    ;    //    sltu x29 x8 x27      ====        sltu t4, s0, s11
                                                  30'd    3535    : data = 32'h    93A16837    ;    //    lui x16 604694      ====        lui a6, 604694
                                                  30'd    3536    : data = 32'h    00BDE933    ;    //    or x18 x27 x11      ====        or s2, s11, a1
                                                  30'd    3537    : data = 32'h    00685933    ;    //    srl x18 x16 x6      ====        srl s2, a6, t1
                                                  30'd    3538    : data = 32'h    40CD5593    ;    //    srai x11 x26 12      ====        srai a1, s10, 12
                                                  30'd    3539    : data = 32'h    ECE6EA13    ;    //    ori x20 x13 -306      ====        ori s4, a3, -306
                                                  30'd    3540    : data = 32'h    01035833    ;    //    srl x16 x6 x16      ====        srl a6, t1, a6
                                                  30'd    3541    : data = 32'h    4064D9B3    ;    //    sra x19 x9 x6      ====        sra s3, s1, t1
                                                  30'd    3542    : data = 32'h    0132BFB3    ;    //    sltu x31 x5 x19      ====        sltu t6, t0, s3
                                                  30'd    3543    : data = 32'h    000DADB3    ;    //    slt x27 x27 x0      ====        slt s11, s11, zero
                                                  30'd    3544    : data = 32'h    EED53E13    ;    //    sltiu x28 x10 -275      ====        sltiu t3, a0, -275
                                                  30'd    3545    : data = 32'h    01A1E633    ;    //    or x12 x3 x26      ====        or a2, gp, s10
                                                  30'd    3546    : data = 32'h    34811937    ;    //    lui x18 215057      ====        lui s2, 215057
                                                  30'd    3547    : data = 32'h    0130A3B3    ;    //    slt x7 x1 x19      ====        slt t2, ra, s3
                                                  30'd    3548    : data = 32'h    49DBC417    ;    //    auipc x8 302524      ====        auipc s0, 302524
                                                  30'd    3549    : data = 32'h    008F8333    ;    //    add x6 x31 x8      ====        add t1, t6, s0
                                                  30'd    3550    : data = 32'h    009741B3    ;    //    xor x3 x14 x9      ====        xor gp, a4, s1
                                                  30'd    3551    : data = 32'h    F4874FB7    ;    //    lui x31 1001588      ====        lui t6, 1001588
                                                  30'd    3552    : data = 32'h    003F2CB3    ;    //    slt x25 x30 x3      ====        slt s9, t5, gp
                                                  30'd    3553    : data = 32'h    012DAE33    ;    //    slt x28 x27 x18      ====        slt t3, s11, s2
                                                  30'd    3554    : data = 32'h    0001E033    ;    //    or x0 x3 x0      ====        or zero, gp, zero
                                                  30'd    3555    : data = 32'h    016DAD33    ;    //    slt x26 x27 x22      ====        slt s10, s11, s6
                                                  30'd    3556    : data = 32'h    F7306B13    ;    //    ori x22 x0 -141      ====        ori s6, zero, -141
                                                  30'd    3557    : data = 32'h    004A8D33    ;    //    add x26 x21 x4      ====        add s10, s5, tp
                                                  30'd    3558    : data = 32'h    85214913    ;    //    xori x18 x2 -1966      ====        xori s2, sp, -1966
                                                  30'd    3559    : data = 32'h    00FDD2B3    ;    //    srl x5 x27 x15      ====        srl t0, s11, a5
                                                  30'd    3560    : data = 32'h    A91CFA13    ;    //    andi x20 x25 -1391      ====        andi s4, s9, -1391
                                                  30'd    3561    : data = 32'h    F65C7D13    ;    //    andi x26 x24 -155      ====        andi s10, s8, -155
                                                  30'd    3562    : data = 32'h    00443433    ;    //    sltu x8 x8 x4      ====        sltu s0, s0, tp
                                                  30'd    3563    : data = 32'h    00D684B3    ;    //    add x9 x13 x13      ====        add s1, a3, a3
                                                  30'd    3564    : data = 32'h    6745A093    ;    //    slti x1 x11 1652      ====        slti ra, a1, 1652
                                                  30'd    3565    : data = 32'h    0C1ECC93    ;    //    xori x25 x29 193      ====        xori s9, t4, 193
                                                  30'd    3566    : data = 32'h    BEF1A113    ;    //    slti x2 x3 -1041      ====        slti sp, gp, -1041
                                                  30'd    3567    : data = 32'h    004D57B3    ;    //    srl x15 x26 x4      ====        srl a5, s10, tp
                                                  30'd    3568    : data = 32'h    379B5817    ;    //    auipc x16 227765      ====        auipc a6, 227765
                                                  30'd    3569    : data = 32'h    0190EFB3    ;    //    or x31 x1 x25      ====        or t6, ra, s9
                                                  30'd    3570    : data = 32'h    01091313    ;    //    slli x6 x18 16      ====        slli t1, s2, 16
                                                  30'd    3571    : data = 32'h    3740A713    ;    //    slti x14 x1 884      ====        slti a4, ra, 884
                                                  30'd    3572    : data = 32'h    EE71BE37    ;    //    lui x28 976667      ====        lui t3, 976667
                                                  30'd    3573    : data = 32'h    000538B3    ;    //    sltu x17 x10 x0      ====        sltu a7, a0, zero
                                                  30'd    3574    : data = 32'h    00526A33    ;    //    or x20 x4 x5      ====        or s4, tp, t0
                                                  30'd    3575    : data = 32'h    417B5D93    ;    //    srai x27 x22 23      ====        srai s11, s6, 23
                                                  30'd    3576    : data = 32'h    01A4FCB3    ;    //    and x25 x9 x26      ====        and s9, s1, s10
                                                  30'd    3577    : data = 32'h    01729913    ;    //    slli x18 x5 23      ====        slli s2, t0, 23
                                                  30'd    3578    : data = 32'h    709969B7    ;    //    lui x19 461206      ====        lui s3, 461206
                                                  30'd    3579    : data = 32'h    41928E33    ;    //    sub x28 x5 x25      ====        sub t3, t0, s9
                                                  30'd    3580    : data = 32'h    78614A17    ;    //    auipc x20 493076      ====        auipc s4, 493076
                                                  30'd    3581    : data = 32'h    DC1C0E97    ;    //    auipc x29 901568      ====        auipc t4, 901568
                                                  30'd    3582    : data = 32'h    402D5693    ;    //    srai x13 x26 2      ====        srai a3, s10, 2
                                                  30'd    3583    : data = 32'h    61D3CB93    ;    //    xori x23 x7 1565      ====        xori s7, t2, 1565
                                                  30'd    3584    : data = 32'h    01BF2933    ;    //    slt x18 x30 x27      ====        slt s2, t5, s11
                                                  30'd    3585    : data = 32'h    A6EC6E37    ;    //    lui x28 683718      ====        lui t3, 683718
                                                  30'd    3586    : data = 32'h    2F716593    ;    //    ori x11 x2 759      ====        ori a1, sp, 759
                                                  30'd    3587    : data = 32'h    30D4E093    ;    //    ori x1 x9 781      ====        ori ra, s1, 781
                                                  30'd    3588    : data = 32'h    00FC9933    ;    //    sll x18 x25 x15      ====        sll s2, s9, a5
                                                  30'd    3589    : data = 32'h    00ADA1B3    ;    //    slt x3 x27 x10      ====        slt gp, s11, a0
                                                  30'd    3590    : data = 32'h    00DC4B33    ;    //    xor x22 x24 x13      ====        xor s6, s8, a3
                                                  30'd    3591    : data = 32'h    3A70AC93    ;    //    slti x25 x1 935      ====        slti s9, ra, 935
                                                  30'd    3592    : data = 32'h    00708833    ;    //    add x16 x1 x7      ====        add a6, ra, t2
                                                  30'd    3593    : data = 32'h    01EDC9B3    ;    //    xor x19 x27 x30      ====        xor s3, s11, t5
                                                  30'd    3594    : data = 32'h    FAFF2713    ;    //    slti x14 x30 -81      ====        slti a4, t5, -81
                                                  30'd    3595    : data = 32'h    41D6D293    ;    //    srai x5 x13 29      ====        srai t0, a3, 29
                                                  30'd    3596    : data = 32'h    8D120C37    ;    //    lui x24 577824      ====        lui s8, 577824
                                                  30'd    3597    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3598    : data = 32'h    00365413    ;    //    srli x8 x12 3      ====        srli s0, a2, 3
                                                  30'd    3599    : data = 32'h    01E2FD33    ;    //    and x26 x5 x30      ====        and s10, t0, t5
                                                  30'd    3600    : data = 32'h    01C283B3    ;    //    add x7 x5 x28      ====        add t2, t0, t3
                                                  30'd    3601    : data = 32'h    00C0DF93    ;    //    srli x31 x1 12      ====        srli t6, ra, 12
                                                  30'd    3602    : data = 32'h    005D7AB3    ;    //    and x21 x26 x5      ====        and s5, s10, t0
                                                  30'd    3603    : data = 32'h    A2CEC293    ;    //    xori x5 x29 -1492      ====        xori t0, t4, -1492
                                                  30'd    3604    : data = 32'h    E4F68913    ;    //    addi x18 x13 -433      ====        addi s2, a3, -433
                                                  30'd    3605    : data = 32'h    0080A2B3    ;    //    slt x5 x1 x8      ====        slt t0, ra, s0
                                                  30'd    3606    : data = 32'h    A04D2793    ;    //    slti x15 x26 -1532      ====        slti a5, s10, -1532
                                                  30'd    3607    : data = 32'h    4184D293    ;    //    srai x5 x9 24      ====        srai t0, s1, 24
                                                  30'd    3608    : data = 32'h    012D1993    ;    //    slli x19 x26 18      ====        slli s3, s10, 18
                                                  30'd    3609    : data = 32'h    00524633    ;    //    xor x12 x4 x5      ====        xor a2, tp, t0
                                                  30'd    3610    : data = 32'h    016FA733    ;    //    slt x14 x31 x22      ====        slt a4, t6, s6
                                                  30'd    3611    : data = 32'h    80000737    ;    //    lui x14 524288      ====        li a4, 0x80000000 #start riscv_int_numeric_corner_stream_17
                                                  30'd    3612    : data = 32'h    00070713    ;    //    addi x14 x14 0      ====        li a4, 0x80000000 #start riscv_int_numeric_corner_stream_17
                                                  30'd    3613    : data = 32'h    15236837    ;    //    lui x16 86582      ====        li a6, 0x152366d5
                                                  30'd    3614    : data = 32'h    6D580813    ;    //    addi x16 x16 1749      ====        li a6, 0x152366d5
                                                  30'd    3615    : data = 32'h    80000B37    ;    //    lui x22 524288      ====        li s6, 0x80000000
                                                  30'd    3616    : data = 32'h    000B0B13    ;    //    addi x22 x22 0      ====        li s6, 0x80000000
                                                  30'd    3617    : data = 32'h    FFF00913    ;    //    addi x18 x0 -1      ====        li s2, 0xffffffff
                                                  30'd    3618    : data = 32'h    00000613    ;    //    addi x12 x0 0      ====        li a2, 0x0
                                                  30'd    3619    : data = 32'h    800005B7    ;    //    lui x11 524288      ====        li a1, 0x80000000
                                                  30'd    3620    : data = 32'h    00058593    ;    //    addi x11 x11 0      ====        li a1, 0x80000000
                                                  30'd    3621    : data = 32'h    00000113    ;    //    addi x2 x0 0      ====        li sp, 0x0
                                                  30'd    3622    : data = 32'h    E7B45BB7    ;    //    lui x23 949061      ====        li s7, 0xe7b44ad9
                                                  30'd    3623    : data = 32'h    AD9B8B93    ;    //    addi x23 x23 -1319      ====        li s7, 0xe7b44ad9
                                                  30'd    3624    : data = 32'h    00000F93    ;    //    addi x31 x0 0      ====        li t6, 0x0
                                                  30'd    3625    : data = 32'h    F49BB7B7    ;    //    lui x15 1001915      ====        li a5, 0xf49bb641
                                                  30'd    3626    : data = 32'h    64178793    ;    //    addi x15 x15 1601      ====        li a5, 0xf49bb641
                                                  30'd    3627    : data = 32'h    A456E837    ;    //    lui x16 673134      ====        lui a6, 673134
                                                  30'd    3628    : data = 32'h    6B270913    ;    //    addi x18 x14 1714      ====        addi s2, a4, 1714
                                                  30'd    3629    : data = 32'h    01F78833    ;    //    add x16 x15 x31      ====        add a6, a5, t6
                                                  30'd    3630    : data = 32'h    412585B3    ;    //    sub x11 x11 x18      ====        sub a1, a1, s2
                                                  30'd    3631    : data = 32'h    7DBC8617    ;    //    auipc x12 515016      ====        auipc a2, 515016
                                                  30'd    3632    : data = 32'h    41F105B3    ;    //    sub x11 x2 x31      ====        sub a1, sp, t6
                                                  30'd    3633    : data = 32'h    63D58593    ;    //    addi x11 x11 1597      ====        addi a1, a1, 1597
                                                  30'd    3634    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3635    : data = 32'h    01F60833    ;    //    add x16 x12 x31      ====        add a6, a2, t6
                                                  30'd    3636    : data = 32'h    C411A837    ;    //    lui x16 803098      ====        lui a6, 803098
                                                  30'd    3637    : data = 32'h    F1DFB817    ;    //    auipc x16 990715      ====        auipc a6, 990715
                                                  30'd    3638    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3639    : data = 32'h    4D710793    ;    //    addi x15 x2 1239      ====        addi a5, sp, 1239
                                                  30'd    3640    : data = 32'h    41780833    ;    //    sub x16 x16 x23      ====        sub a6, a6, s7
                                                  30'd    3641    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3642    : data = 32'h    00F90633    ;    //    add x12 x18 x15      ====        add a2, s2, a5
                                                  30'd    3643    : data = 32'h    412F8633    ;    //    sub x12 x31 x18      ====        sub a2, t6, s2
                                                  30'd    3644    : data = 32'h    41FB8133    ;    //    sub x2 x23 x31      ====        sub sp, s7, t6
                                                  30'd    3645    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3646    : data = 32'h    0B832FB7    ;    //    lui x31 47154      ====        lui t6, 47154
                                                  30'd    3647    : data = 32'h    01080BB3    ;    //    add x23 x16 x16      ====        add s7, a6, a6
                                                  30'd    3648    : data = 32'h    CB1F8793    ;    //    addi x15 x31 -847      ====        addi a5, t6, -847
                                                  30'd    3649    : data = 32'h    18C01617    ;    //    auipc x12 101377      ====        auipc a2, 101377
                                                  30'd    3650    : data = 32'h    40B80933    ;    //    sub x18 x16 x11      ====        sub s2, a6, a1
                                                  30'd    3651    : data = 32'h    41F907B3    ;    //    sub x15 x18 x31      ====        sub a5, s2, t6
                                                  30'd    3652    : data = 32'h    317F8813    ;    //    addi x16 x31 791      ====        addi a6, t6, 791
                                                  30'd    3653    : data = 32'h    4B690793    ;    //    addi x15 x18 1206      ====        addi a5, s2, 1206
                                                  30'd    3654    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3655    : data = 32'h    5CD070EF    ;    //    jal x1 32204      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_17
                                                  30'd    3656    : data = 32'h    61A86593    ;    //    ori x11 x16 1562      ====        ori a1, a6, 1562
                                                  30'd    3657    : data = 32'h    48598B13    ;    //    addi x22 x19 1157      ====        addi s6, s3, 1157
                                                  30'd    3658    : data = 32'h    01990D33    ;    //    add x26 x18 x25      ====        add s10, s2, s9
                                                  30'd    3659    : data = 32'h    001C51B3    ;    //    srl x3 x24 x1      ====        srl gp, s8, ra
                                                  30'd    3660    : data = 32'h    2D6DEA93    ;    //    ori x21 x27 726      ====        ori s5, s11, 726
                                                  30'd    3661    : data = 32'h    41400733    ;    //    sub x14 x0 x20      ====        sub a4, zero, s4
                                                  30'd    3662    : data = 32'h    41DADDB3    ;    //    sra x27 x21 x29      ====        sra s11, s5, t4
                                                  30'd    3663    : data = 32'h    7DE8BD93    ;    //    sltiu x27 x17 2014      ====        sltiu s11, a7, 2014
                                                  30'd    3664    : data = 32'h    20DFD337    ;    //    lui x6 134653      ====        lui t1, 134653
                                                  30'd    3665    : data = 32'h    41F651B3    ;    //    sra x3 x12 x31      ====        sra gp, a2, t6
                                                  30'd    3666    : data = 32'h    58A20B93    ;    //    addi x23 x4 1418      ====        addi s7, tp, 1418
                                                  30'd    3667    : data = 32'h    87908BB7    ;    //    lui x23 555272      ====        lui s7, 555272
                                                  30'd    3668    : data = 32'h    CFBFBC93    ;    //    sltiu x25 x31 -773      ====        sltiu s9, t6, -773
                                                  30'd    3669    : data = 32'h    4184D913    ;    //    srai x18 x9 24      ====        srai s2, s1, 24
                                                  30'd    3670    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3671    : data = 32'h    4025D913    ;    //    srai x18 x11 2      ====        srai s2, a1, 2
                                                  30'd    3672    : data = 32'h    01307D33    ;    //    and x26 x0 x19      ====        and s10, zero, s3
                                                  30'd    3673    : data = 32'h    411E5493    ;    //    srai x9 x28 17      ====        srai s1, t3, 17
                                                  30'd    3674    : data = 32'h    004FDDB3    ;    //    srl x27 x31 x4      ====        srl s11, t6, tp
                                                  30'd    3675    : data = 32'h    A23B6A97    ;    //    auipc x21 664502      ====        auipc s5, 664502
                                                  30'd    3676    : data = 32'h    001178B3    ;    //    and x17 x2 x1      ====        and a7, sp, ra
                                                  30'd    3677    : data = 32'h    003FD5B3    ;    //    srl x11 x31 x3      ====        srl a1, t6, gp
                                                  30'd    3678    : data = 32'h    017DAD33    ;    //    slt x26 x27 x23      ====        slt s10, s11, s7
                                                  30'd    3679    : data = 32'h    C9513897    ;    //    auipc x17 824595      ====        auipc a7, 824595
                                                  30'd    3680    : data = 32'h    77176197    ;    //    auipc x3 487798      ====        auipc gp, 487798
                                                  30'd    3681    : data = 32'h    AF76A313    ;    //    slti x6 x13 -1289      ====        slti t1, a3, -1289
                                                  30'd    3682    : data = 32'h    7855E797    ;    //    auipc x15 492894      ====        auipc a5, 492894
                                                  30'd    3683    : data = 32'h    00385713    ;    //    srli x14 x16 3      ====        srli a4, a6, 3
                                                  30'd    3684    : data = 32'h    01A6EB33    ;    //    or x22 x13 x26      ====        or s6, a3, s10
                                                  30'd    3685    : data = 32'h    00180833    ;    //    add x16 x16 x1      ====        add a6, a6, ra
                                                  30'd    3686    : data = 32'h    9946A993    ;    //    slti x19 x13 -1644      ====        slti s3, a3, -1644
                                                  30'd    3687    : data = 32'h    0183D133    ;    //    srl x2 x7 x24      ====        srl sp, t2, s8
                                                  30'd    3688    : data = 32'h    0A08BC93    ;    //    sltiu x25 x17 160      ====        sltiu s9, a7, 160
                                                  30'd    3689    : data = 32'h    01D52B33    ;    //    slt x22 x10 x29      ====        slt s6, a0, t4
                                                  30'd    3690    : data = 32'h    D53DE193    ;    //    ori x3 x27 -685      ====        ori gp, s11, -685
                                                  30'd    3691    : data = 32'h    7147A493    ;    //    slti x9 x15 1812      ====        slti s1, a5, 1812
                                                  30'd    3692    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3693    : data = 32'h    00D4DB13    ;    //    srli x22 x9 13      ====        srli s6, s1, 13
                                                  30'd    3694    : data = 32'h    40E8D813    ;    //    srai x16 x17 14      ====        srai a6, a7, 14
                                                  30'd    3695    : data = 32'h    F3564037    ;    //    lui x0 996708      ====        lui zero, 996708
                                                  30'd    3696    : data = 32'h    00427AB3    ;    //    and x21 x4 x4      ====        and s5, tp, tp
                                                  30'd    3697    : data = 32'h    01C6DB13    ;    //    srli x22 x13 28      ====        srli s6, a3, 28
                                                  30'd    3698    : data = 32'h    E8FDFE13    ;    //    andi x28 x27 -369      ====        andi t3, s11, -369
                                                  30'd    3699    : data = 32'h    E3F06113    ;    //    ori x2 x0 -449      ====        ori sp, zero, -449
                                                  30'd    3700    : data = 32'h    01AB4733    ;    //    xor x14 x22 x26      ====        xor a4, s6, s10
                                                  30'd    3701    : data = 32'h    418DD2B3    ;    //    sra x5 x27 x24      ====        sra t0, s11, s8
                                                  30'd    3702    : data = 32'h    008921B3    ;    //    slt x3 x18 x8      ====        slt gp, s2, s0
                                                  30'd    3703    : data = 32'h    9A342D13    ;    //    slti x26 x8 -1629      ====        slti s10, s0, -1629
                                                  30'd    3704    : data = 32'h    01F96133    ;    //    or x2 x18 x31      ====        or sp, s2, t6
                                                  30'd    3705    : data = 32'h    ADE7B393    ;    //    sltiu x7 x15 -1314      ====        sltiu t2, a5, -1314
                                                  30'd    3706    : data = 32'h    01230EB3    ;    //    add x29 x6 x18      ====        add t4, t1, s2
                                                  30'd    3707    : data = 32'h    0083D093    ;    //    srli x1 x7 8      ====        srli ra, t2, 8
                                                  30'd    3708    : data = 32'h    4012D893    ;    //    srai x17 x5 1      ====        srai a7, t0, 1
                                                  30'd    3709    : data = 32'h    00EEFA33    ;    //    and x20 x29 x14      ====        and s4, t4, a4
                                                  30'd    3710    : data = 32'h    0045F3B3    ;    //    and x7 x11 x4      ====        and t2, a1, tp
                                                  30'd    3711    : data = 32'h    0199CD33    ;    //    xor x26 x19 x25      ====        xor s10, s3, s9
                                                  30'd    3712    : data = 32'h    01AE74B3    ;    //    and x9 x28 x26      ====        and s1, t3, s10
                                                  30'd    3713    : data = 32'h    7B892DB7    ;    //    lui x27 506002      ====        lui s11, 506002
                                                  30'd    3714    : data = 32'h    018F99B3    ;    //    sll x19 x31 x24      ====        sll s3, t6, s8
                                                  30'd    3715    : data = 32'h    01ACCDB3    ;    //    xor x27 x25 x26      ====        xor s11, s9, s10
                                                  30'd    3716    : data = 32'h    40DA8CB3    ;    //    sub x25 x21 x13      ====        sub s9, s5, a3
                                                  30'd    3717    : data = 32'h    A0F74B13    ;    //    xori x22 x14 -1521      ====        xori s6, a4, -1521
                                                  30'd    3718    : data = 32'h    8F05C493    ;    //    xori x9 x11 -1808      ====        xori s1, a1, -1808
                                                  30'd    3719    : data = 32'h    2E7AF393    ;    //    andi x7 x21 743      ====        andi t2, s5, 743
                                                  30'd    3720    : data = 32'h    00D5CC33    ;    //    xor x24 x11 x13      ====        xor s8, a1, a3
                                                  30'd    3721    : data = 32'h    15F6FDB7    ;    //    lui x27 89967      ====        lui s11, 89967
                                                  30'd    3722    : data = 32'h    00AF52B3    ;    //    srl x5 x30 x10      ====        srl t0, t5, a0
                                                  30'd    3723    : data = 32'h    473AE413    ;    //    ori x8 x21 1139      ====        ori s0, s5, 1139
                                                  30'd    3724    : data = 32'h    A96F0C13    ;    //    addi x24 x30 -1386      ====        addi s8, t5, -1386
                                                  30'd    3725    : data = 32'h    00195D93    ;    //    srli x27 x18 1      ====        srli s11, s2, 1
                                                  30'd    3726    : data = 32'h    0082B833    ;    //    sltu x16 x5 x8      ====        sltu a6, t0, s0
                                                  30'd    3727    : data = 32'h    68BF7013    ;    //    andi x0 x30 1675      ====        andi zero, t5, 1675
                                                  30'd    3728    : data = 32'h    011A5933    ;    //    srl x18 x20 x17      ====        srl s2, s4, a7
                                                  30'd    3729    : data = 32'h    00161033    ;    //    sll x0 x12 x1      ====        sll zero, a2, ra
                                                  30'd    3730    : data = 32'h    40B680B3    ;    //    sub x1 x13 x11      ====        sub ra, a3, a1
                                                  30'd    3731    : data = 32'h    5F68D337    ;    //    lui x6 390797      ====        lui t1, 390797
                                                  30'd    3732    : data = 32'h    409ED2B3    ;    //    sra x5 x29 x9      ====        sra t0, t4, s1
                                                  30'd    3733    : data = 32'h    00346A33    ;    //    or x20 x8 x3      ====        or s4, s0, gp
                                                  30'd    3734    : data = 32'h    01981C13    ;    //    slli x24 x16 25      ====        slli s8, a6, 25
                                                  30'd    3735    : data = 32'h    01E64733    ;    //    xor x14 x12 x30      ====        xor a4, a2, t5
                                                  30'd    3736    : data = 32'h    0016A433    ;    //    slt x8 x13 x1      ====        slt s0, a3, ra
                                                  30'd    3737    : data = 32'h    01DDA033    ;    //    slt x0 x27 x29      ====        slt zero, s11, t4
                                                  30'd    3738    : data = 32'h    55E14613    ;    //    xori x12 x2 1374      ====        xori a2, sp, 1374
                                                  30'd    3739    : data = 32'h    76ABCA13    ;    //    xori x20 x23 1898      ====        xori s4, s7, 1898
                                                  30'd    3740    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3741    : data = 32'h    012F0333    ;    //    add x6 x30 x18      ====        add t1, t5, s2
                                                  30'd    3742    : data = 32'h    0100FE33    ;    //    and x28 x1 x16      ====        and t3, ra, a6
                                                  30'd    3743    : data = 32'h    01D62633    ;    //    slt x12 x12 x29      ====        slt a2, a2, t4
                                                  30'd    3744    : data = 32'h    0125B1B3    ;    //    sltu x3 x11 x18      ====        sltu gp, a1, s2
                                                  30'd    3745    : data = 32'h    B9784C13    ;    //    xori x24 x16 -1129      ====        xori s8, a6, -1129
                                                  30'd    3746    : data = 32'h    C1C50293    ;    //    addi x5 x10 -996      ====        addi t0, a0, -996
                                                  30'd    3747    : data = 32'h    120224B7    ;    //    lui x9 73762      ====        lui s1, 73762
                                                  30'd    3748    : data = 32'h    01795733    ;    //    srl x14 x18 x23      ====        srl a4, s2, s7
                                                  30'd    3749    : data = 32'h    B7DC0C13    ;    //    addi x24 x24 -1155      ====        addi s8, s8, -1155
                                                  30'd    3750    : data = 32'h    52D18C37    ;    //    lui x24 339224      ====        lui s8, 339224
                                                  30'd    3751    : data = 32'h    96464C13    ;    //    xori x24 x12 -1692      ====        xori s8, a2, -1692
                                                  30'd    3752    : data = 32'h    01F51BB3    ;    //    sll x23 x10 x31      ====        sll s7, a0, t6
                                                  30'd    3753    : data = 32'h    407A03B3    ;    //    sub x7 x20 x7      ====        sub t2, s4, t2
                                                  30'd    3754    : data = 32'h    00C29713    ;    //    slli x14 x5 12      ====        slli a4, t0, 12
                                                  30'd    3755    : data = 32'h    0157B033    ;    //    sltu x0 x15 x21      ====        sltu zero, a5, s5
                                                  30'd    3756    : data = 32'h    D1979297    ;    //    auipc x5 858489      ====        auipc t0, 858489
                                                  30'd    3757    : data = 32'h    01D728B3    ;    //    slt x17 x14 x29      ====        slt a7, a4, t4
                                                  30'd    3758    : data = 32'h    F04B4493    ;    //    xori x9 x22 -252      ====        xori s1, s6, -252
                                                  30'd    3759    : data = 32'h    E513BD93    ;    //    sltiu x27 x7 -431      ====        sltiu s11, t2, -431
                                                  30'd    3760    : data = 32'h    00CF32B3    ;    //    sltu x5 x30 x12      ====        sltu t0, t5, a2
                                                  30'd    3761    : data = 32'h    D37ED6B7    ;    //    lui x13 866285      ====        lui a3, 866285
                                                  30'd    3762    : data = 32'h    0E8D4413    ;    //    xori x8 x26 232      ====        xori s0, s10, 232
                                                  30'd    3763    : data = 32'h    F3BD0693    ;    //    addi x13 x26 -197      ====        addi a3, s10, -197
                                                  30'd    3764    : data = 32'h    00D91193    ;    //    slli x3 x18 13      ====        slli gp, s2, 13
                                                  30'd    3765    : data = 32'h    40D15913    ;    //    srai x18 x2 13      ====        srai s2, sp, 13
                                                  30'd    3766    : data = 32'h    01F6B833    ;    //    sltu x16 x13 x31      ====        sltu a6, a3, t6
                                                  30'd    3767    : data = 32'h    008AA0B3    ;    //    slt x1 x21 x8      ====        slt ra, s5, s0
                                                  30'd    3768    : data = 32'h    004217B3    ;    //    sll x15 x4 x4      ====        sll a5, tp, tp
                                                  30'd    3769    : data = 32'h    005D0833    ;    //    add x16 x26 x5      ====        add a6, s10, t0
                                                  30'd    3770    : data = 32'h    60449B37    ;    //    lui x22 394313      ====        lui s6, 394313
                                                  30'd    3771    : data = 32'h    003F1A13    ;    //    slli x20 x30 3      ====        slli s4, t5, 3
                                                  30'd    3772    : data = 32'h    005A1293    ;    //    slli x5 x20 5      ====        slli t0, s4, 5
                                                  30'd    3773    : data = 32'h    0131D6B3    ;    //    srl x13 x3 x19      ====        srl a3, gp, s3
                                                  30'd    3774    : data = 32'h    01EB6833    ;    //    or x16 x22 x30      ====        or a6, s6, t5
                                                  30'd    3775    : data = 32'h    4113D7B3    ;    //    sra x15 x7 x17      ====        sra a5, t2, a7
                                                  30'd    3776    : data = 32'h    41BA5BB3    ;    //    sra x23 x20 x27      ====        sra s7, s4, s11
                                                  30'd    3777    : data = 32'h    7C54AB13    ;    //    slti x22 x9 1989      ====        slti s6, s1, 1989
                                                  30'd    3778    : data = 32'h    00002933    ;    //    slt x18 x0 x0      ====        slt s2, zero, zero
                                                  30'd    3779    : data = 32'h    EB842F93    ;    //    slti x31 x8 -328      ====        slti t6, s0, -328
                                                  30'd    3780    : data = 32'h    00F605B3    ;    //    add x11 x12 x15      ====        add a1, a2, a5
                                                  30'd    3781    : data = 32'h    5EB08913    ;    //    addi x18 x1 1515      ====        addi s2, ra, 1515
                                                  30'd    3782    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3783    : data = 32'h    00C8C2B3    ;    //    xor x5 x17 x12      ====        xor t0, a7, a2
                                                  30'd    3784    : data = 32'h    A88F3E37    ;    //    lui x28 690419      ====        lui t3, 690419
                                                  30'd    3785    : data = 32'h    4024D913    ;    //    srai x18 x9 2      ====        srai s2, s1, 2
                                                  30'd    3786    : data = 32'h    01BC5833    ;    //    srl x16 x24 x27      ====        srl a6, s8, s11
                                                  30'd    3787    : data = 32'h    44732497    ;    //    auipc x9 280370      ====        auipc s1, 280370
                                                  30'd    3788    : data = 32'h    28EAE713    ;    //    ori x14 x21 654      ====        ori a4, s5, 654
                                                  30'd    3789    : data = 32'h    006B9093    ;    //    slli x1 x23 6      ====        slli ra, s7, 6
                                                  30'd    3790    : data = 32'h    00765EB3    ;    //    srl x29 x12 x7      ====        srl t4, a2, t2
                                                  30'd    3791    : data = 32'h    01A09113    ;    //    slli x2 x1 26      ====        slli sp, ra, 26
                                                  30'd    3792    : data = 32'h    80000B37    ;    //    lui x22 524288      ====        li s6, 0x80000000 #start riscv_int_numeric_corner_stream_34
                                                  30'd    3793    : data = 32'h    000B0B13    ;    //    addi x22 x22 0      ====        li s6, 0x80000000 #start riscv_int_numeric_corner_stream_34
                                                  30'd    3794    : data = 32'h    E51DBC37    ;    //    lui x24 938459      ====        li s8, 0xe51dae1e
                                                  30'd    3795    : data = 32'h    E1EC0C13    ;    //    addi x24 x24 -482      ====        li s8, 0xe51dae1e
                                                  30'd    3796    : data = 32'h    00000393    ;    //    addi x7 x0 0      ====        li t2, 0x0
                                                  30'd    3797    : data = 32'h    00000593    ;    //    addi x11 x0 0      ====        li a1, 0x0
                                                  30'd    3798    : data = 32'h    FFF00E93    ;    //    addi x29 x0 -1      ====        li t4, 0xffffffff
                                                  30'd    3799    : data = 32'h    FFF00493    ;    //    addi x9 x0 -1      ====        li s1, 0xffffffff
                                                  30'd    3800    : data = 32'h    58588A37    ;    //    lui x20 361864      ====        li s4, 0x58588507
                                                  30'd    3801    : data = 32'h    507A0A13    ;    //    addi x20 x20 1287      ====        li s4, 0x58588507
                                                  30'd    3802    : data = 32'h    00000793    ;    //    addi x15 x0 0      ====        li a5, 0x0
                                                  30'd    3803    : data = 32'h    00000E13    ;    //    addi x28 x0 0      ====        li t3, 0x0
                                                  30'd    3804    : data = 32'h    00000613    ;    //    addi x12 x0 0      ====        li a2, 0x0
                                                  30'd    3805    : data = 32'h    8C4E8793    ;    //    addi x15 x29 -1852      ====        addi a5, t4, -1852
                                                  30'd    3806    : data = 32'h    BD3B0C13    ;    //    addi x24 x22 -1069      ====        addi s8, s6, -1069
                                                  30'd    3807    : data = 32'h    12F0D637    ;    //    lui x12 77581      ====        lui a2, 77581
                                                  30'd    3808    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3809    : data = 32'h    F8658613    ;    //    addi x12 x11 -122      ====        addi a2, a1, -122
                                                  30'd    3810    : data = 32'h    C9D26C17    ;    //    auipc x24 826662      ====        auipc s8, 826662
                                                  30'd    3811    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3812    : data = 32'h    01CE84B3    ;    //    add x9 x29 x28      ====        add s1, t4, t3
                                                  30'd    3813    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3814    : data = 32'h    007B0A33    ;    //    add x20 x22 x7      ====        add s4, s6, t2
                                                  30'd    3815    : data = 32'h    A88CE797    ;    //    auipc x15 690382      ====        auipc a5, 690382
                                                  30'd    3816    : data = 32'h    01C583B3    ;    //    add x7 x11 x28      ====        add t2, a1, t3
                                                  30'd    3817    : data = 32'h    40F583B3    ;    //    sub x7 x11 x15      ====        sub t2, a1, a5
                                                  30'd    3818    : data = 32'h    9AA0FC17    ;    //    auipc x24 633359      ====        auipc s8, 633359
                                                  30'd    3819    : data = 32'h    416385B3    ;    //    sub x11 x7 x22      ====        sub a1, t2, s6
                                                  30'd    3820    : data = 32'h    016783B3    ;    //    add x7 x15 x22      ====        add t2, a5, s6
                                                  30'd    3821    : data = 32'h    AEE7E3B7    ;    //    lui x7 716414      ====        lui t2, 716414
                                                  30'd    3822    : data = 32'h    00938B33    ;    //    add x22 x7 x9      ====        add s6, t2, s1
                                                  30'd    3823    : data = 32'h    32D070EF    ;    //    jal x1 31532      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_34
                                                  30'd    3824    : data = 32'h    003F7B33    ;    //    and x22 x30 x3      ====        and s6, t5, gp
                                                  30'd    3825    : data = 32'h    6FC58A13    ;    //    addi x20 x11 1788      ====        addi s4, a1, 1788
                                                  30'd    3826    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3827    : data = 32'h    00EADFB3    ;    //    srl x31 x21 x14      ====        srl t6, s5, a4
                                                  30'd    3828    : data = 32'h    01232B33    ;    //    slt x22 x6 x18      ====        slt s6, t1, s2
                                                  30'd    3829    : data = 32'h    C5947A37    ;    //    lui x20 809287      ====        lui s4, 809287
                                                  30'd    3830    : data = 32'h    40CB5B13    ;    //    srai x22 x22 12      ====        srai s6, s6, 12
                                                  30'd    3831    : data = 32'h    01B60DB3    ;    //    add x27 x12 x27      ====        add s11, a2, s11
                                                  30'd    3832    : data = 32'h    01E21113    ;    //    slli x2 x4 30      ====        slli sp, tp, 30
                                                  30'd    3833    : data = 32'h    01B3D133    ;    //    srl x2 x7 x27      ====        srl sp, t2, s11
                                                  30'd    3834    : data = 32'h    00757CB3    ;    //    and x25 x10 x7      ====        and s9, a0, t2
                                                  30'd    3835    : data = 32'h    01E68833    ;    //    add x16 x13 x30      ====        add a6, a3, t5
                                                  30'd    3836    : data = 32'h    598A4F93    ;    //    xori x31 x20 1432      ====        xori t6, s4, 1432
                                                  30'd    3837    : data = 32'h    40C452B3    ;    //    sra x5 x8 x12      ====        sra t0, s0, a2
                                                  30'd    3838    : data = 32'h    4099DF93    ;    //    srai x31 x19 9      ====        srai t6, s3, 9
                                                  30'd    3839    : data = 32'h    00785113    ;    //    srli x2 x16 7      ====        srli sp, a6, 7
                                                  30'd    3840    : data = 32'h    4183D893    ;    //    srai x17 x7 24      ====        srai a7, t2, 24
                                                  30'd    3841    : data = 32'h    B3EB0713    ;    //    addi x14 x22 -1218      ====        addi a4, s6, -1218
                                                  30'd    3842    : data = 32'h    1BC27313    ;    //    andi x6 x4 444      ====        andi t1, tp, 444
                                                  30'd    3843    : data = 32'h    BA674B93    ;    //    xori x23 x14 -1114      ====        xori s7, a4, -1114
                                                  30'd    3844    : data = 32'h    006CD5B3    ;    //    srl x11 x25 x6      ====        srl a1, s9, t1
                                                  30'd    3845    : data = 32'h    00B70333    ;    //    add x6 x14 x11      ====        add t1, a4, a1
                                                  30'd    3846    : data = 32'h    0026A333    ;    //    slt x6 x13 x2      ====        slt t1, a3, sp
                                                  30'd    3847    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3848    : data = 32'h    0113E733    ;    //    or x14 x7 x17      ====        or a4, t2, a7
                                                  30'd    3849    : data = 32'h    00D56DB3    ;    //    or x27 x10 x13      ====        or s11, a0, a3
                                                  30'd    3850    : data = 32'h    00CB8DB3    ;    //    add x27 x23 x12      ====        add s11, s7, a2
                                                  30'd    3851    : data = 32'h    14623393    ;    //    sltiu x7 x4 326      ====        sltiu t2, tp, 326
                                                  30'd    3852    : data = 32'h    71F72B17    ;    //    auipc x22 466802      ====        auipc s6, 466802
                                                  30'd    3853    : data = 32'h    00EE4933    ;    //    xor x18 x28 x14      ====        xor s2, t3, a4
                                                  30'd    3854    : data = 32'h    011D9913    ;    //    slli x18 x27 17      ====        slli s2, s11, 17
                                                  30'd    3855    : data = 32'h    007A58B3    ;    //    srl x17 x20 x7      ====        srl a7, s4, t2
                                                  30'd    3856    : data = 32'h    005446B3    ;    //    xor x13 x8 x5      ====        xor a3, s0, t0
                                                  30'd    3857    : data = 32'h    38E4E293    ;    //    ori x5 x9 910      ====        ori t0, s1, 910
                                                  30'd    3858    : data = 32'h    F2DB3113    ;    //    sltiu x2 x22 -211      ====        sltiu sp, s6, -211
                                                  30'd    3859    : data = 32'h    081BC913    ;    //    xori x18 x23 129      ====        xori s2, s7, 129
                                                  30'd    3860    : data = 32'h    D9607E93    ;    //    andi x29 x0 -618      ====        andi t4, zero, -618
                                                  30'd    3861    : data = 32'h    0114C133    ;    //    xor x2 x9 x17      ====        xor sp, s1, a7
                                                  30'd    3862    : data = 32'h    00399B93    ;    //    slli x23 x19 3      ====        slli s7, s3, 3
                                                  30'd    3863    : data = 32'h    4C757D13    ;    //    andi x26 x10 1223      ====        andi s10, a0, 1223
                                                  30'd    3864    : data = 32'h    01DF36B3    ;    //    sltu x13 x30 x29      ====        sltu a3, t5, t4
                                                  30'd    3865    : data = 32'h    017772B3    ;    //    and x5 x14 x23      ====        and t0, a4, s7
                                                  30'd    3866    : data = 32'h    007F4333    ;    //    xor x6 x30 x7      ====        xor t1, t5, t2
                                                  30'd    3867    : data = 32'h    00E74933    ;    //    xor x18 x14 x14      ====        xor s2, a4, a4
                                                  30'd    3868    : data = 32'h    41FCD593    ;    //    srai x11 x25 31      ====        srai a1, s9, 31
                                                  30'd    3869    : data = 32'h    01C9E3B3    ;    //    or x7 x19 x28      ====        or t2, s3, t3
                                                  30'd    3870    : data = 32'h    0044B433    ;    //    sltu x8 x9 x4      ====        sltu s0, s1, tp
                                                  30'd    3871    : data = 32'h    009C7C33    ;    //    and x24 x24 x9      ====        and s8, s8, s1
                                                  30'd    3872    : data = 32'h    1D954193    ;    //    xori x3 x10 473      ====        xori gp, a0, 473
                                                  30'd    3873    : data = 32'h    000776B3    ;    //    and x13 x14 x0      ====        and a3, a4, zero
                                                  30'd    3874    : data = 32'h    41C8D2B3    ;    //    sra x5 x17 x28      ====        sra t0, a7, t3
                                                  30'd    3875    : data = 32'h    00981D33    ;    //    sll x26 x16 x9      ====        sll s10, a6, s1
                                                  30'd    3876    : data = 32'h    00115F93    ;    //    srli x31 x2 1      ====        srli t6, sp, 1
                                                  30'd    3877    : data = 32'h    00829D13    ;    //    slli x26 x5 8      ====        slli s10, t0, 8
                                                  30'd    3878    : data = 32'h    005C8133    ;    //    add x2 x25 x5      ====        add sp, s9, t0
                                                  30'd    3879    : data = 32'h    00E69A93    ;    //    slli x21 x13 14      ====        slli s5, a3, 14
                                                  30'd    3880    : data = 32'h    406B5C93    ;    //    srai x25 x22 6      ====        srai s9, s6, 6
                                                  30'd    3881    : data = 32'h    403B0E33    ;    //    sub x28 x22 x3      ====        sub t3, s6, gp
                                                  30'd    3882    : data = 32'h    23BA7E13    ;    //    andi x28 x20 571      ====        andi t3, s4, 571
                                                  30'd    3883    : data = 32'h    29407493    ;    //    andi x9 x0 660      ====        andi s1, zero, 660
                                                  30'd    3884    : data = 32'h    0149AAB3    ;    //    slt x21 x19 x20      ====        slt s5, s3, s4
                                                  30'd    3885    : data = 32'h    9042B417    ;    //    auipc x8 590891      ====        auipc s0, 590891
                                                  30'd    3886    : data = 32'h    84097413    ;    //    andi x8 x18 -1984      ====        andi s0, s2, -1984
                                                  30'd    3887    : data = 32'h    003BC1B3    ;    //    xor x3 x23 x3      ====        xor gp, s7, gp
                                                  30'd    3888    : data = 32'h    01AC33B3    ;    //    sltu x7 x24 x26      ====        sltu t2, s8, s10
                                                  30'd    3889    : data = 32'h    40400CB3    ;    //    sub x25 x0 x4      ====        sub s9, zero, tp
                                                  30'd    3890    : data = 32'h    01535713    ;    //    srli x14 x6 21      ====        srli a4, t1, 21
                                                  30'd    3891    : data = 32'h    AE1A4C13    ;    //    xori x24 x20 -1311      ====        xori s8, s4, -1311
                                                  30'd    3892    : data = 32'h    00E1D933    ;    //    srl x18 x3 x14      ====        srl s2, gp, a4
                                                  30'd    3893    : data = 32'h    4067D633    ;    //    sra x12 x15 x6      ====        sra a2, a5, t1
                                                  30'd    3894    : data = 32'h    496A0B93    ;    //    addi x23 x20 1174      ====        addi s7, s4, 1174
                                                  30'd    3895    : data = 32'h    013A42B3    ;    //    xor x5 x20 x19      ====        xor t0, s4, s3
                                                  30'd    3896    : data = 32'h    40E55413    ;    //    srai x8 x10 14      ====        srai s0, a0, 14
                                                  30'd    3897    : data = 32'h    D9484313    ;    //    xori x6 x16 -620      ====        xori t1, a6, -620
                                                  30'd    3898    : data = 32'h    D2663C93    ;    //    sltiu x25 x12 -730      ====        sltiu s9, a2, -730
                                                  30'd    3899    : data = 32'h    857AC993    ;    //    xori x19 x21 -1961      ====        xori s3, s5, -1961
                                                  30'd    3900    : data = 32'h    005FE1B3    ;    //    or x3 x31 x5      ====        or gp, t6, t0
                                                  30'd    3901    : data = 32'h    0171CA33    ;    //    xor x20 x3 x23      ====        xor s4, gp, s7
                                                  30'd    3902    : data = 32'h    41EDD033    ;    //    sra x0 x27 x30      ====        sra zero, s11, t5
                                                  30'd    3903    : data = 32'h    0036ADB3    ;    //    slt x27 x13 x3      ====        slt s11, a3, gp
                                                  30'd    3904    : data = 32'h    00927433    ;    //    and x8 x4 x9      ====        and s0, tp, s1
                                                  30'd    3905    : data = 32'h    9DE6A293    ;    //    slti x5 x13 -1570      ====        slti t0, a3, -1570
                                                  30'd    3906    : data = 32'h    FE610293    ;    //    addi x5 x2 -26      ====        addi t0, sp, -26
                                                  30'd    3907    : data = 32'h    000D4B33    ;    //    xor x22 x26 x0      ====        xor s6, s10, zero
                                                  30'd    3908    : data = 32'h    418E5033    ;    //    sra x0 x28 x24      ====        sra zero, t3, s8
                                                  30'd    3909    : data = 32'h    01B19593    ;    //    slli x11 x3 27      ====        slli a1, gp, 27
                                                  30'd    3910    : data = 32'h    0174DF93    ;    //    srli x31 x9 23      ====        srli t6, s1, 23
                                                  30'd    3911    : data = 32'h    00442633    ;    //    slt x12 x8 x4      ====        slt a2, s0, tp
                                                  30'd    3912    : data = 32'h    01B4E8B3    ;    //    or x17 x9 x27      ====        or a7, s1, s11
                                                  30'd    3913    : data = 32'h    C0872E37    ;    //    lui x28 788594      ====        lui t3, 788594
                                                  30'd    3914    : data = 32'h    00990733    ;    //    add x14 x18 x9      ====        add a4, s2, s1
                                                  30'd    3915    : data = 32'h    C19DE293    ;    //    ori x5 x27 -999      ====        ori t0, s11, -999
                                                  30'd    3916    : data = 32'h    8EE4F793    ;    //    andi x15 x9 -1810      ====        andi a5, s1, -1810
                                                  30'd    3917    : data = 32'h    4089DCB3    ;    //    sra x25 x19 x8      ====        sra s9, s3, s0
                                                  30'd    3918    : data = 32'h    86D4E693    ;    //    ori x13 x9 -1939      ====        ori a3, s1, -1939
                                                  30'd    3919    : data = 32'h    2FFA2B93    ;    //    slti x23 x20 767      ====        slti s7, s4, 767
                                                  30'd    3920    : data = 32'h    00CB5333    ;    //    srl x6 x22 x12      ====        srl t1, s6, a2
                                                  30'd    3921    : data = 32'h    360E6D13    ;    //    ori x26 x28 864      ====        ori s10, t3, 864
                                                  30'd    3922    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3923    : data = 32'h    FE894893    ;    //    xori x17 x18 -24      ====        xori a7, s2, -24
                                                  30'd    3924    : data = 32'h    AC79BE97    ;    //    auipc x29 706459      ====        auipc t4, 706459
                                                  30'd    3925    : data = 32'h    157A0A13    ;    //    addi x20 x20 343      ====        addi s4, s4, 343
                                                  30'd    3926    : data = 32'h    00725093    ;    //    srli x1 x4 7      ====        srli ra, tp, 7
                                                  30'd    3927    : data = 32'h    64329337    ;    //    lui x6 410409      ====        lui t1, 410409
                                                  30'd    3928    : data = 32'h    407E0B33    ;    //    sub x22 x28 x7      ====        sub s6, t3, t2
                                                  30'd    3929    : data = 32'h    41760AB3    ;    //    sub x21 x12 x23      ====        sub s5, a2, s7
                                                  30'd    3930    : data = 32'h    5DBEBC93    ;    //    sltiu x25 x29 1499      ====        sltiu s9, t4, 1499
                                                  30'd    3931    : data = 32'h    5856FE93    ;    //    andi x29 x13 1413      ====        andi t4, a3, 1413
                                                  30'd    3932    : data = 32'h    1FBC6913    ;    //    ori x18 x24 507      ====        ori s2, s8, 507
                                                  30'd    3933    : data = 32'h    CFC31937    ;    //    lui x18 850993      ====        lui s2, 850993
                                                  30'd    3934    : data = 32'h    08090393    ;    //    addi x7 x18 128      ====        addi t2, s2, 128
                                                  30'd    3935    : data = 32'h    40C9D433    ;    //    sra x8 x19 x12      ====        sra s0, s3, a2
                                                  30'd    3936    : data = 32'h    F7F11DB7    ;    //    lui x27 1015569      ====        lui s11, 1015569
                                                  30'd    3937    : data = 32'h    C3AAEE93    ;    //    ori x29 x21 -966      ====        ori t4, s5, -966
                                                  30'd    3938    : data = 32'h    84637E13    ;    //    andi x28 x6 -1978      ====        andi t3, t1, -1978
                                                  30'd    3939    : data = 32'h    41040B33    ;    //    sub x22 x8 x16      ====        sub s6, s0, a6
                                                  30'd    3940    : data = 32'h    9DBAD3B7    ;    //    lui x7 646061      ====        lui t2, 646061
                                                  30'd    3941    : data = 32'h    019FF2B3    ;    //    and x5 x31 x25      ====        and t0, t6, s9
                                                  30'd    3942    : data = 32'h    00B05F93    ;    //    srli x31 x0 11      ====        srli t6, zero, 11
                                                  30'd    3943    : data = 32'h    98C78C93    ;    //    addi x25 x15 -1652      ====        addi s9, a5, -1652
                                                  30'd    3944    : data = 32'h    0067F0B3    ;    //    and x1 x15 x6      ====        and ra, a5, t1
                                                  30'd    3945    : data = 32'h    F05AAC13    ;    //    slti x24 x21 -251      ====        slti s8, s5, -251
                                                  30'd    3946    : data = 32'h    0FB14093    ;    //    xori x1 x2 251      ====        xori ra, sp, 251
                                                  30'd    3947    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3948    : data = 32'h    35743D93    ;    //    sltiu x27 x8 855      ====        sltiu s11, s0, 855
                                                  30'd    3949    : data = 32'h    7BDAA593    ;    //    slti x11 x21 1981      ====        slti a1, s5, 1981
                                                  30'd    3950    : data = 32'h    0007A333    ;    //    slt x6 x15 x0      ====        slt t1, a5, zero
                                                  30'd    3951    : data = 32'h    00FA5A13    ;    //    srli x20 x20 15      ====        srli s4, s4, 15
                                                  30'd    3952    : data = 32'h    FAA5FC17    ;    //    auipc x24 1026655      ====        auipc s8, 1026655
                                                  30'd    3953    : data = 32'h    0FA5B713    ;    //    sltiu x14 x11 250      ====        sltiu a4, a1, 250
                                                  30'd    3954    : data = 32'h    40818EB3    ;    //    sub x29 x3 x8      ====        sub t4, gp, s0
                                                  30'd    3955    : data = 32'h    01C583B3    ;    //    add x7 x11 x28      ====        add t2, a1, t3
                                                  30'd    3956    : data = 32'h    01681D33    ;    //    sll x26 x16 x22      ====        sll s10, a6, s6
                                                  30'd    3957    : data = 32'h    018E2BB3    ;    //    slt x23 x28 x24      ====        slt s7, t3, s8
                                                  30'd    3958    : data = 32'h    415E5313    ;    //    srai x6 x28 21      ====        srai t1, t3, 21
                                                  30'd    3959    : data = 32'h    00D5EAB3    ;    //    or x21 x11 x13      ====        or s5, a1, a3
                                                  30'd    3960    : data = 32'h    652ABE93    ;    //    sltiu x29 x21 1618      ====        sltiu t4, s5, 1618
                                                  30'd    3961    : data = 32'h    7306AE17    ;    //    auipc x28 471146      ====        auipc t3, 471146
                                                  30'd    3962    : data = 32'h    006089B3    ;    //    add x19 x1 x6      ====        add s3, ra, t1
                                                  30'd    3963    : data = 32'h    8B850793    ;    //    addi x15 x10 -1864      ====        addi a5, a0, -1864
                                                  30'd    3964    : data = 32'h    0137F133    ;    //    and x2 x15 x19      ====        and sp, a5, s3
                                                  30'd    3965    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3966    : data = 32'h    41F80933    ;    //    sub x18 x16 x31      ====        sub s2, a6, t6
                                                  30'd    3967    : data = 32'h    01760933    ;    //    add x18 x12 x23      ====        add s2, a2, s7
                                                  30'd    3968    : data = 32'h    032EA613    ;    //    slti x12 x29 50      ====        slti a2, t4, 50
                                                  30'd    3969    : data = 32'h    D7BB4397    ;    //    auipc x7 883636      ====        auipc t2, 883636
                                                  30'd    3970    : data = 32'h    81D14793    ;    //    xori x15 x2 -2019      ====        xori a5, sp, -2019
                                                  30'd    3971    : data = 32'h    71DDFE17    ;    //    auipc x28 466399      ====        auipc t3, 466399
                                                  30'd    3972    : data = 32'h    F76C4893    ;    //    xori x17 x24 -138      ====        xori a7, s8, -138
                                                  30'd    3973    : data = 32'h    D1D0A837    ;    //    lui x16 859402      ====        lui a6, 859402
                                                  30'd    3974    : data = 32'h    0134EEB3    ;    //    or x29 x9 x19      ====        or t4, s1, s3
                                                  30'd    3975    : data = 32'h    D5DA7017    ;    //    auipc x0 875943      ====        auipc zero, 875943
                                                  30'd    3976    : data = 32'h    017E92B3    ;    //    sll x5 x29 x23      ====        sll t0, t4, s7
                                                  30'd    3977    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    3978    : data = 32'h    CD230993    ;    //    addi x19 x6 -814      ====        addi s3, t1, -814
                                                  30'd    3979    : data = 32'h    00AC1393    ;    //    slli x7 x24 10      ====        slli t2, s8, 10
                                                  30'd    3980    : data = 32'h    018ED713    ;    //    srli x14 x29 24      ====        srli a4, t4, 24
                                                  30'd    3981    : data = 32'h    36D6B717    ;    //    auipc x14 224619      ====        auipc a4, 224619
                                                  30'd    3982    : data = 32'h    EFDECCB7    ;    //    lui x25 982508      ====        lui s9, 982508
                                                  30'd    3983    : data = 32'h    01595013    ;    //    srli x0 x18 21      ====        srli zero, s2, 21
                                                  30'd    3984    : data = 32'h    A3F8C813    ;    //    xori x16 x17 -1473      ====        xori a6, a7, -1473
                                                  30'd    3985    : data = 32'h    405B8AB3    ;    //    sub x21 x23 x5      ====        sub s5, s7, t0
                                                  30'd    3986    : data = 32'h    01A35933    ;    //    srl x18 x6 x26      ====        srl s2, t1, s10
                                                  30'd    3987    : data = 32'h    EE35E317    ;    //    auipc x6 975710      ====        auipc t1, 975710
                                                  30'd    3988    : data = 32'h    40568D33    ;    //    sub x26 x13 x5      ====        sub s10, a3, t0
                                                  30'd    3989    : data = 32'h    68A9DD37    ;    //    lui x26 428701      ====        lui s10, 428701
                                                  30'd    3990    : data = 32'h    6000A593    ;    //    slti x11 x1 1536      ====        slti a1, ra, 1536
                                                  30'd    3991    : data = 32'h    008AA8B3    ;    //    slt x17 x21 x8      ====        slt a7, s5, s0
                                                  30'd    3992    : data = 32'h    1500A613    ;    //    slti x12 x1 336      ====        slti a2, ra, 336
                                                  30'd    3993    : data = 32'h    0CA3FD93    ;    //    andi x27 x7 202      ====        andi s11, t2, 202
                                                  30'd    3994    : data = 32'h    BACBBD13    ;    //    sltiu x26 x23 -1108      ====        sltiu s10, s7, -1108
                                                  30'd    3995    : data = 32'h    40A75813    ;    //    srai x16 x14 10      ====        srai a6, a4, 10
                                                  30'd    3996    : data = 32'h    C26A4593    ;    //    xori x11 x20 -986      ====        xori a1, s4, -986
                                                  30'd    3997    : data = 32'h    41EC84B3    ;    //    sub x9 x25 x30      ====        sub s1, s9, t5
                                                  30'd    3998    : data = 32'h    416A8E33    ;    //    sub x28 x21 x22      ====        sub t3, s5, s6
                                                  30'd    3999    : data = 32'h    01C185B3    ;    //    add x11 x3 x28      ====        add a1, gp, t3
                                                  30'd    4000    : data = 32'h    7BDBC893    ;    //    xori x17 x23 1981      ====        xori a7, s7, 1981
                                                  30'd    4001    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4002    : data = 32'h    11FD4113    ;    //    xori x2 x26 287      ====        xori sp, s10, 287
                                                  30'd    4003    : data = 32'h    A1EC37B7    ;    //    lui x15 663235      ====        lui a5, 663235
                                                  30'd    4004    : data = 32'h    01CEECB3    ;    //    or x25 x29 x28      ====        or s9, t4, t3
                                                  30'd    4005    : data = 32'h    48733D93    ;    //    sltiu x27 x6 1159      ====        sltiu s11, t1, 1159
                                                  30'd    4006    : data = 32'h    003E6C33    ;    //    or x24 x28 x3      ====        or s8, t3, gp
                                                  30'd    4007    : data = 32'h    41715633    ;    //    sra x12 x2 x23      ====        sra a2, sp, s7
                                                  30'd    4008    : data = 32'h    3A48C613    ;    //    xori x12 x17 932      ====        xori a2, a7, 932
                                                  30'd    4009    : data = 32'h    01C50EB3    ;    //    add x29 x10 x28      ====        add t4, a0, t3
                                                  30'd    4010    : data = 32'h    27BDC613    ;    //    xori x12 x27 635      ====        xori a2, s11, 635
                                                  30'd    4011    : data = 32'h    5E49F713    ;    //    andi x14 x19 1508      ====        andi a4, s3, 1508
                                                  30'd    4012    : data = 32'h    00EA44B3    ;    //    xor x9 x20 x14      ====        xor s1, s4, a4
                                                  30'd    4013    : data = 32'h    00C5D193    ;    //    srli x3 x11 12      ====        srli gp, a1, 12
                                                  30'd    4014    : data = 32'h    002E5833    ;    //    srl x16 x28 x2      ====        srl a6, t3, sp
                                                  30'd    4015    : data = 32'h    01178033    ;    //    add x0 x15 x17      ====        add zero, a5, a7
                                                  30'd    4016    : data = 32'h    1E3F0613    ;    //    addi x12 x30 483      ====        addi a2, t5, 483
                                                  30'd    4017    : data = 32'h    01857DB3    ;    //    and x27 x10 x24      ====        and s11, a0, s8
                                                  30'd    4018    : data = 32'h    01F674B3    ;    //    and x9 x12 x31      ====        and s1, a2, t6
                                                  30'd    4019    : data = 32'h    8E5A2893    ;    //    slti x17 x20 -1819      ====        slti a7, s4, -1819
                                                  30'd    4020    : data = 32'h    0F60C713    ;    //    xori x14 x1 246      ====        xori a4, ra, 246
                                                  30'd    4021    : data = 32'h    25AE4397    ;    //    auipc x7 154340      ====        auipc t2, 154340
                                                  30'd    4022    : data = 32'h    FDDDCC13    ;    //    xori x24 x27 -35      ====        xori s8, s11, -35
                                                  30'd    4023    : data = 32'h    00CC0E33    ;    //    add x28 x24 x12      ====        add t3, s8, a2
                                                  30'd    4024    : data = 32'h    6067AB13    ;    //    slti x22 x15 1542      ====        slti s6, a5, 1542
                                                  30'd    4025    : data = 32'h    01094FB3    ;    //    xor x31 x18 x16      ====        xor t6, s2, a6
                                                  30'd    4026    : data = 32'h    0538B813    ;    //    sltiu x16 x17 83      ====        sltiu a6, a7, 83
                                                  30'd    4027    : data = 32'h    00025E93    ;    //    srli x29 x4 0      ====        srli t4, tp, 0
                                                  30'd    4028    : data = 32'h    40C15913    ;    //    srai x18 x2 12      ====        srai s2, sp, 12
                                                  30'd    4029    : data = 32'h    01341733    ;    //    sll x14 x8 x19      ====        sll a4, s0, s3
                                                  30'd    4030    : data = 32'h    008277B3    ;    //    and x15 x4 x8      ====        and a5, tp, s0
                                                  30'd    4031    : data = 32'h    00FB53B3    ;    //    srl x7 x22 x15      ====        srl t2, s6, a5
                                                  30'd    4032    : data = 32'h    C4ECAD93    ;    //    slti x27 x25 -946      ====        slti s11, s9, -946
                                                  30'd    4033    : data = 32'h    3415B613    ;    //    sltiu x12 x11 833      ====        sltiu a2, a1, 833
                                                  30'd    4034    : data = 32'h    00559993    ;    //    slli x19 x11 5      ====        slli s3, a1, 5
                                                  30'd    4035    : data = 32'h    92AEA093    ;    //    slti x1 x29 -1750      ====        slti ra, t4, -1750
                                                  30'd    4036    : data = 32'h    00CD55B3    ;    //    srl x11 x26 x12      ====        srl a1, s10, a2
                                                  30'd    4037    : data = 32'h    30EEEA97    ;    //    auipc x21 200430      ====        auipc s5, 200430
                                                  30'd    4038    : data = 32'h    00037833    ;    //    and x16 x6 x0      ====        and a6, t1, zero
                                                  30'd    4039    : data = 32'h    019A5133    ;    //    srl x2 x20 x25      ====        srl sp, s4, s9
                                                  30'd    4040    : data = 32'h    03E16393    ;    //    ori x7 x2 62      ====        ori t2, sp, 62
                                                  30'd    4041    : data = 32'h    01FD8433    ;    //    add x8 x27 x31      ====        add s0, s11, t6
                                                  30'd    4042    : data = 32'h    B8D10A93    ;    //    addi x21 x2 -1139      ====        addi s5, sp, -1139
                                                  30'd    4043    : data = 32'h    00F24FB3    ;    //    xor x31 x4 x15      ====        xor t6, tp, a5
                                                  30'd    4044    : data = 32'h    413453B3    ;    //    sra x7 x8 x19      ====        sra t2, s0, s3
                                                  30'd    4045    : data = 32'h    D9A23117    ;    //    auipc x2 891427      ====        auipc sp, 891427
                                                  30'd    4046    : data = 32'h    013BC7B3    ;    //    xor x15 x23 x19      ====        xor a5, s7, s3
                                                  30'd    4047    : data = 32'h    00FAB833    ;    //    sltu x16 x21 x15      ====        sltu a6, s5, a5
                                                  30'd    4048    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4049    : data = 32'h    94E68313    ;    //    addi x6 x13 -1714      ====        addi t1, a3, -1714
                                                  30'd    4050    : data = 32'h    9E159717    ;    //    auipc x14 647513      ====        auipc a4, 647513
                                                  30'd    4051    : data = 32'h    00F668B3    ;    //    or x17 x12 x15      ====        or a7, a2, a5
                                                  30'd    4052    : data = 32'h    2B120037    ;    //    lui x0 176416      ====        lui zero, 176416
                                                  30'd    4053    : data = 32'h    431A0893    ;    //    addi x17 x20 1073      ====        addi a7, s4, 1073
                                                  30'd    4054    : data = 32'h    DEB2A113    ;    //    slti x2 x5 -533      ====        slti sp, t0, -533
                                                  30'd    4055    : data = 32'h    AB32C817    ;    //    auipc x16 701228      ====        auipc a6, 701228
                                                  30'd    4056    : data = 32'h    016CA8B3    ;    //    slt x17 x25 x22      ====        slt a7, s9, s6
                                                  30'd    4057    : data = 32'h    E9348593    ;    //    addi x11 x9 -365      ====        addi a1, s1, -365
                                                  30'd    4058    : data = 32'h    5893CE93    ;    //    xori x29 x7 1417      ====        xori t4, t2, 1417
                                                  30'd    4059    : data = 32'h    010196B3    ;    //    sll x13 x3 x16      ====        sll a3, gp, a6
                                                  30'd    4060    : data = 32'h    01F46033    ;    //    or x0 x8 x31      ====        or zero, s0, t6
                                                  30'd    4061    : data = 32'h    DE5FF313    ;    //    andi x6 x31 -539      ====        andi t1, t6, -539
                                                  30'd    4062    : data = 32'h    9D55E093    ;    //    ori x1 x11 -1579      ====        ori ra, a1, -1579
                                                  30'd    4063    : data = 32'h    A7D73293    ;    //    sltiu x5 x14 -1411      ====        sltiu t0, a4, -1411
                                                  30'd    4064    : data = 32'h    AA58CB17    ;    //    auipc x22 697740      ====        auipc s6, 697740
                                                  30'd    4065    : data = 32'h    41BE8433    ;    //    sub x8 x29 x27      ====        sub s0, t4, s11
                                                  30'd    4066    : data = 32'h    01AC1633    ;    //    sll x12 x24 x26      ====        sll a2, s8, s10
                                                  30'd    4067    : data = 32'h    01C1FC33    ;    //    and x24 x3 x28      ====        and s8, gp, t3
                                                  30'd    4068    : data = 32'h    01066DB3    ;    //    or x27 x12 x16      ====        or s11, a2, a6
                                                  30'd    4069    : data = 32'h    00EF9B13    ;    //    slli x22 x31 14      ====        slli s6, t6, 14
                                                  30'd    4070    : data = 32'h    002AFEB3    ;    //    and x29 x21 x2      ====        and t4, s5, sp
                                                  30'd    4071    : data = 32'h    EDF82C93    ;    //    slti x25 x16 -289      ====        slti s9, a6, -289
                                                  30'd    4072    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4073    : data = 32'h    41F75813    ;    //    srai x16 x14 31      ====        srai a6, a4, 31
                                                  30'd    4074    : data = 32'h    409457B3    ;    //    sra x15 x8 x9      ====        sra a5, s0, s1
                                                  30'd    4075    : data = 32'h    414E02B3    ;    //    sub x5 x28 x20      ====        sub t0, t3, s4
                                                  30'd    4076    : data = 32'h    8E2EFB37    ;    //    lui x22 582383      ====        lui s6, 582383
                                                  30'd    4077    : data = 32'h    886F8593    ;    //    addi x11 x31 -1914      ====        addi a1, t6, -1914
                                                  30'd    4078    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4079    : data = 32'h    2C5AEB13    ;    //    ori x22 x21 709      ====        ori s6, s5, 709
                                                  30'd    4080    : data = 32'h    418DDE13    ;    //    srai x28 x27 24      ====        srai t3, s11, 24
                                                  30'd    4081    : data = 32'h    00005193    ;    //    srli x3 x0 0      ====        srli gp, zero, 0
                                                  30'd    4082    : data = 32'h    79A8A813    ;    //    slti x16 x17 1946      ====        slti a6, a7, 1946
                                                  30'd    4083    : data = 32'h    B7768713    ;    //    addi x14 x13 -1161      ====        addi a4, a3, -1161
                                                  30'd    4084    : data = 32'h    008F9D93    ;    //    slli x27 x31 8      ====        slli s11, t6, 8
                                                  30'd    4085    : data = 32'h    41C25B33    ;    //    sra x22 x4 x28      ====        sra s6, tp, t3
                                                  30'd    4086    : data = 32'h    410C88B3    ;    //    sub x17 x25 x16      ====        sub a7, s9, a6
                                                  30'd    4087    : data = 32'h    6E940B93    ;    //    addi x23 x8 1769      ====        addi s7, s0, 1769
                                                  30'd    4088    : data = 32'h    012F5033    ;    //    srl x0 x30 x18      ====        srl zero, t5, s2
                                                  30'd    4089    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4090    : data = 32'h    00B68833    ;    //    add x16 x13 x11      ====        add a6, a3, a1
                                                  30'd    4091    : data = 32'h    01B08B33    ;    //    add x22 x1 x27      ====        add s6, ra, s11
                                                  30'd    4092    : data = 32'h    4969A293    ;    //    slti x5 x19 1174      ====        slti t0, s3, 1174
                                                  30'd    4093    : data = 32'h    81B93D13    ;    //    sltiu x26 x18 -2021      ====        sltiu s10, s2, -2021
                                                  30'd    4094    : data = 32'h    00AA7B33    ;    //    and x22 x20 x10      ====        and s6, s4, a0
                                                  30'd    4095    : data = 32'h    CFF7E593    ;    //    ori x11 x15 -769      ====        ori a1, a5, -769
                                                  30'd    4096    : data = 32'h    41D25A93    ;    //    srai x21 x4 29      ====        srai s5, tp, 29
                                                  30'd    4097    : data = 32'h    015A80B3    ;    //    add x1 x21 x21      ====        add ra, s5, s5
                                                  30'd    4098    : data = 32'h    0008D9B3    ;    //    srl x19 x17 x0      ====        srl s3, a7, zero
                                                  30'd    4099    : data = 32'h    54208C13    ;    //    addi x24 x1 1346      ====        addi s8, ra, 1346
                                                  30'd    4100    : data = 32'h    1D42AE13    ;    //    slti x28 x5 468      ====        slti t3, t0, 468
                                                  30'd    4101    : data = 32'h    0145EEB3    ;    //    or x29 x11 x20      ====        or t4, a1, s4
                                                  30'd    4102    : data = 32'h    008F63B3    ;    //    or x7 x30 x8      ====        or t2, t5, s0
                                                  30'd    4103    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4104    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4105    : data = 32'h    6774A293    ;    //    slti x5 x9 1655      ====        slti t0, s1, 1655
                                                  30'd    4106    : data = 32'h    40DF59B3    ;    //    sra x19 x30 x13      ====        sra s3, t5, a3
                                                  30'd    4107    : data = 32'h    01721B13    ;    //    slli x22 x4 23      ====        slli s6, tp, 23
                                                  30'd    4108    : data = 32'h    010309B3    ;    //    add x19 x6 x16      ====        add s3, t1, a6
                                                  30'd    4109    : data = 32'h    01FC0333    ;    //    add x6 x24 x31      ====        add t1, s8, t6
                                                  30'd    4110    : data = 32'h    004552B3    ;    //    srl x5 x10 x4      ====        srl t0, a0, tp
                                                  30'd    4111    : data = 32'h    E7BA0113    ;    //    addi x2 x20 -389      ====        addi sp, s4, -389
                                                  30'd    4112    : data = 32'h    A7884093    ;    //    xori x1 x16 -1416      ====        xori ra, a6, -1416
                                                  30'd    4113    : data = 32'h    0097B633    ;    //    sltu x12 x15 x9      ====        sltu a2, a5, s1
                                                  30'd    4114    : data = 32'h    01FD5333    ;    //    srl x6 x26 x31      ====        srl t1, s10, t6
                                                  30'd    4115    : data = 32'h    BA2EC117    ;    //    auipc x2 762604      ====        auipc sp, 762604
                                                  30'd    4116    : data = 32'h    80000737    ;    //    lui x14 524288      ====        li a4, 0x80000000 #start riscv_int_numeric_corner_stream_18
                                                  30'd    4117    : data = 32'h    00070713    ;    //    addi x14 x14 0      ====        li a4, 0x80000000 #start riscv_int_numeric_corner_stream_18
                                                  30'd    4118    : data = 32'h    1491D6B7    ;    //    lui x13 84253      ====        li a3, 0x1491c988
                                                  30'd    4119    : data = 32'h    98868693    ;    //    addi x13 x13 -1656      ====        li a3, 0x1491c988
                                                  30'd    4120    : data = 32'h    00000D93    ;    //    addi x27 x0 0      ====        li s11, 0x0
                                                  30'd    4121    : data = 32'h    80000CB7    ;    //    lui x25 524288      ====        li s9, 0x80000000
                                                  30'd    4122    : data = 32'h    000C8C93    ;    //    addi x25 x25 0      ====        li s9, 0x80000000
                                                  30'd    4123    : data = 32'h    00000A13    ;    //    addi x20 x0 0      ====        li s4, 0x0
                                                  30'd    4124    : data = 32'h    00000413    ;    //    addi x8 x0 0      ====        li s0, 0x0
                                                  30'd    4125    : data = 32'h    00000C13    ;    //    addi x24 x0 0      ====        li s8, 0x0
                                                  30'd    4126    : data = 32'h    FFF00293    ;    //    addi x5 x0 -1      ====        li t0, 0xffffffff
                                                  30'd    4127    : data = 32'h    FA702137    ;    //    lui x2 1025794      ====        li sp, 0xfa701cfd
                                                  30'd    4128    : data = 32'h    CFD10113    ;    //    addi x2 x2 -771      ====        li sp, 0xfa701cfd
                                                  30'd    4129    : data = 32'h    3146F837    ;    //    lui x16 201839      ====        li a6, 0x3146ef54
                                                  30'd    4130    : data = 32'h    F5480813    ;    //    addi x16 x16 -172      ====        li a6, 0x3146ef54
                                                  30'd    4131    : data = 32'h    35008A37    ;    //    lui x20 217096      ====        lui s4, 217096
                                                  30'd    4132    : data = 32'h    92C80D97    ;    //    auipc x27 601216      ====        auipc s11, 601216
                                                  30'd    4133    : data = 32'h    DBEF8817    ;    //    auipc x16 900856      ====        auipc a6, 900856
                                                  30'd    4134    : data = 32'h    2E267CB7    ;    //    lui x25 189031      ====        lui s9, 189031
                                                  30'd    4135    : data = 32'h    290C9A37    ;    //    lui x20 168137      ====        lui s4, 168137
                                                  30'd    4136    : data = 32'h    01940833    ;    //    add x16 x8 x25      ====        add a6, s0, s9
                                                  30'd    4137    : data = 32'h    D0A75117    ;    //    auipc x2 854645      ====        auipc sp, 854645
                                                  30'd    4138    : data = 32'h    418406B3    ;    //    sub x13 x8 x24      ====        sub a3, s0, s8
                                                  30'd    4139    : data = 32'h    40580CB3    ;    //    sub x25 x16 x5      ====        sub s9, a6, t0
                                                  30'd    4140    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4141    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4142    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4143    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4144    : data = 32'h    01980433    ;    //    add x8 x16 x25      ====        add s0, a6, s9
                                                  30'd    4145    : data = 32'h    68C8BC37    ;    //    lui x24 429195      ====        lui s8, 429195
                                                  30'd    4146    : data = 32'h    414D82B3    ;    //    sub x5 x27 x20      ====        sub t0, s11, s4
                                                  30'd    4147    : data = 32'h    61C070EF    ;    //    jal x1 30236      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_18
                                                  30'd    4148    : data = 32'h    0094C633    ;    //    xor x12 x9 x9      ====        xor a2, s1, s1
                                                  30'd    4149    : data = 32'h    B83355B7    ;    //    lui x11 754485      ====        lui a1, 754485
                                                  30'd    4150    : data = 32'h    C0850617    ;    //    auipc x12 788560      ====        auipc a2, 788560
                                                  30'd    4151    : data = 32'h    006D9F93    ;    //    slli x31 x27 6      ====        slli t6, s11, 6
                                                  30'd    4152    : data = 32'h    F4F49797    ;    //    auipc x15 1003337      ====        auipc a5, 1003337
                                                  30'd    4153    : data = 32'h    008606B3    ;    //    add x13 x12 x8      ====        add a3, a2, s0
                                                  30'd    4154    : data = 32'h    F2568913    ;    //    addi x18 x13 -219      ====        addi s2, a3, -219
                                                  30'd    4155    : data = 32'h    6D60CA93    ;    //    xori x21 x1 1750      ====        xori s5, ra, 1750
                                                  30'd    4156    : data = 32'h    014361B3    ;    //    or x3 x6 x20      ====        or gp, t1, s4
                                                  30'd    4157    : data = 32'h    016C2CB3    ;    //    slt x25 x24 x22      ====        slt s9, s8, s6
                                                  30'd    4158    : data = 32'h    84B63593    ;    //    sltiu x11 x12 -1973      ====        sltiu a1, a2, -1973
                                                  30'd    4159    : data = 32'h    0063FB33    ;    //    and x22 x7 x6      ====        and s6, t2, t1
                                                  30'd    4160    : data = 32'h    F1D78D93    ;    //    addi x27 x15 -227      ====        addi s11, a5, -227
                                                  30'd    4161    : data = 32'h    012F5833    ;    //    srl x16 x30 x18      ====        srl a6, t5, s2
                                                  30'd    4162    : data = 32'h    40C353B3    ;    //    sra x7 x6 x12      ====        sra t2, t1, a2
                                                  30'd    4163    : data = 32'h    00065C13    ;    //    srli x24 x12 0      ====        srli s8, a2, 0
                                                  30'd    4164    : data = 32'h    411389B3    ;    //    sub x19 x7 x17      ====        sub s3, t2, a7
                                                  30'd    4165    : data = 32'h    01C0F0B3    ;    //    and x1 x1 x28      ====        and ra, ra, t3
                                                  30'd    4166    : data = 32'h    000B9793    ;    //    slli x15 x23 0      ====        slli a5, s7, 0
                                                  30'd    4167    : data = 32'h    00919933    ;    //    sll x18 x3 x9      ====        sll s2, gp, s1
                                                  30'd    4168    : data = 32'h    014D08B3    ;    //    add x17 x26 x20      ====        add a7, s10, s4
                                                  30'd    4169    : data = 32'h    FEB0E293    ;    //    ori x5 x1 -21      ====        ori t0, ra, -21
                                                  30'd    4170    : data = 32'h    0154F033    ;    //    and x0 x9 x21      ====        and zero, s1, s5
                                                  30'd    4171    : data = 32'h    40B95333    ;    //    sra x6 x18 x11      ====        sra t1, s2, a1
                                                  30'd    4172    : data = 32'h    0D598E93    ;    //    addi x29 x19 213      ====        addi t4, s3, 213
                                                  30'd    4173    : data = 32'h    017CFDB3    ;    //    and x27 x25 x23      ====        and s11, s9, s7
                                                  30'd    4174    : data = 32'h    00B3E833    ;    //    or x16 x7 x11      ====        or a6, t2, a1
                                                  30'd    4175    : data = 32'h    00AD8FB3    ;    //    add x31 x27 x10      ====        add t6, s11, a0
                                                  30'd    4176    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4177    : data = 32'h    011B8833    ;    //    add x16 x23 x17      ====        add a6, s7, a7
                                                  30'd    4178    : data = 32'h    00115933    ;    //    srl x18 x2 x1      ====        srl s2, sp, ra
                                                  30'd    4179    : data = 32'h    8D8ECA13    ;    //    xori x20 x29 -1832      ====        xori s4, t4, -1832
                                                  30'd    4180    : data = 32'h    3CA3AC13    ;    //    slti x24 x7 970      ====        slti s8, t2, 970
                                                  30'd    4181    : data = 32'h    01885733    ;    //    srl x14 x16 x24      ====        srl a4, a6, s8
                                                  30'd    4182    : data = 32'h    B30FC093    ;    //    xori x1 x31 -1232      ====        xori ra, t6, -1232
                                                  30'd    4183    : data = 32'h    40EC5593    ;    //    srai x11 x24 14      ====        srai a1, s8, 14
                                                  30'd    4184    : data = 32'h    014E3433    ;    //    sltu x8 x28 x20      ====        sltu s0, t3, s4
                                                  30'd    4185    : data = 32'h    BB090B13    ;    //    addi x22 x18 -1104      ====        addi s6, s2, -1104
                                                  30'd    4186    : data = 32'h    6224B413    ;    //    sltiu x8 x9 1570      ====        sltiu s0, s1, 1570
                                                  30'd    4187    : data = 32'h    0147DDB3    ;    //    srl x27 x15 x20      ====        srl s11, a5, s4
                                                  30'd    4188    : data = 32'h    18023913    ;    //    sltiu x18 x4 384      ====        sltiu s2, tp, 384
                                                  30'd    4189    : data = 32'h    009BCDB3    ;    //    xor x27 x23 x9      ====        xor s11, s7, s1
                                                  30'd    4190    : data = 32'h    01DA5B13    ;    //    srli x22 x20 29      ====        srli s6, s4, 29
                                                  30'd    4191    : data = 32'h    8FD6A893    ;    //    slti x17 x13 -1795      ====        slti a7, a3, -1795
                                                  30'd    4192    : data = 32'h    015B6033    ;    //    or x0 x22 x21      ====        or zero, s6, s5
                                                  30'd    4193    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4194    : data = 32'h    B20E5617    ;    //    auipc x12 729317      ====        auipc a2, 729317
                                                  30'd    4195    : data = 32'h    01F46C33    ;    //    or x24 x8 x31      ====        or s8, s0, t6
                                                  30'd    4196    : data = 32'h    01A6D493    ;    //    srli x9 x13 26      ====        srli s1, a3, 26
                                                  30'd    4197    : data = 32'h    01239593    ;    //    slli x11 x7 18      ====        slli a1, t2, 18
                                                  30'd    4198    : data = 32'h    01F22B33    ;    //    slt x22 x4 x31      ====        slt s6, tp, t6
                                                  30'd    4199    : data = 32'h    4109DA33    ;    //    sra x20 x19 x16      ====        sra s4, s3, a6
                                                  30'd    4200    : data = 32'h    001B5D93    ;    //    srli x27 x22 1      ====        srli s11, s6, 1
                                                  30'd    4201    : data = 32'h    6D340CB7    ;    //    lui x25 447296      ====        lui s9, 447296
                                                  30'd    4202    : data = 32'h    00E54AB3    ;    //    xor x21 x10 x14      ====        xor s5, a0, a4
                                                  30'd    4203    : data = 32'h    00201E13    ;    //    slli x28 x0 2      ====        slli t3, zero, 2
                                                  30'd    4204    : data = 32'h    716BA113    ;    //    slti x2 x23 1814      ====        slti sp, s7, 1814
                                                  30'd    4205    : data = 32'h    E785CD13    ;    //    xori x26 x11 -392      ====        xori s10, a1, -392
                                                  30'd    4206    : data = 32'h    002222B3    ;    //    slt x5 x4 x2      ====        slt t0, tp, sp
                                                  30'd    4207    : data = 32'h    015324B3    ;    //    slt x9 x6 x21      ====        slt s1, t1, s5
                                                  30'd    4208    : data = 32'h    00769B13    ;    //    slli x22 x13 7      ====        slli s6, a3, 7
                                                  30'd    4209    : data = 32'h    A56C3B13    ;    //    sltiu x22 x24 -1450      ====        sltiu s6, s8, -1450
                                                  30'd    4210    : data = 32'h    E0ECE393    ;    //    ori x7 x25 -498      ====        ori t2, s9, -498
                                                  30'd    4211    : data = 32'h    01E80833    ;    //    add x16 x16 x30      ====        add a6, a6, t5
                                                  30'd    4212    : data = 32'h    01A58733    ;    //    add x14 x11 x26      ====        add a4, a1, s10
                                                  30'd    4213    : data = 32'h    57989297    ;    //    auipc x5 358793      ====        auipc t0, 358793
                                                  30'd    4214    : data = 32'h    D2F4D297    ;    //    auipc x5 864077      ====        auipc t0, 864077
                                                  30'd    4215    : data = 32'h    24A4A0B7    ;    //    lui x1 150090      ====        lui ra, 150090
                                                  30'd    4216    : data = 32'h    01B00633    ;    //    add x12 x0 x27      ====        add a2, zero, s11
                                                  30'd    4217    : data = 32'h    2E2ABEB7    ;    //    lui x29 189099      ====        lui t4, 189099
                                                  30'd    4218    : data = 32'h    00EDC5B3    ;    //    xor x11 x27 x14      ====        xor a1, s11, a4
                                                  30'd    4219    : data = 32'h    233CA913    ;    //    slti x18 x25 563      ====        slti s2, s9, 563
                                                  30'd    4220    : data = 32'h    0133E4B3    ;    //    or x9 x7 x19      ====        or s1, t2, s3
                                                  30'd    4221    : data = 32'h    010E5733    ;    //    srl x14 x28 x16      ====        srl a4, t3, a6
                                                  30'd    4222    : data = 32'h    00E11333    ;    //    sll x6 x2 x14      ====        sll t1, sp, a4
                                                  30'd    4223    : data = 32'h    41985433    ;    //    sra x8 x16 x25      ====        sra s0, a6, s9
                                                  30'd    4224    : data = 32'h    41ABDB93    ;    //    srai x23 x23 26      ====        srai s7, s7, 26
                                                  30'd    4225    : data = 32'h    41265133    ;    //    sra x2 x12 x18      ====        sra sp, a2, s2
                                                  30'd    4226    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4227    : data = 32'h    0099EB33    ;    //    or x22 x19 x9      ====        or s6, s3, s1
                                                  30'd    4228    : data = 32'h    018A62B3    ;    //    or x5 x20 x24      ====        or t0, s4, s8
                                                  30'd    4229    : data = 32'h    B46CEE13    ;    //    ori x28 x25 -1210      ====        ori t3, s9, -1210
                                                  30'd    4230    : data = 32'h    013A9133    ;    //    sll x2 x21 x19      ====        sll sp, s5, s3
                                                  30'd    4231    : data = 32'h    003D21B3    ;    //    slt x3 x26 x3      ====        slt gp, s10, gp
                                                  30'd    4232    : data = 32'h    C5FABA93    ;    //    sltiu x21 x21 -929      ====        sltiu s5, s5, -929
                                                  30'd    4233    : data = 32'h    015180B3    ;    //    add x1 x3 x21      ====        add ra, gp, s5
                                                  30'd    4234    : data = 32'h    01509E33    ;    //    sll x28 x1 x21      ====        sll t3, ra, s5
                                                  30'd    4235    : data = 32'h    00C52BB3    ;    //    slt x23 x10 x12      ====        slt s7, a0, a2
                                                  30'd    4236    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4237    : data = 32'h    00C8D113    ;    //    srli x2 x17 12      ====        srli sp, a7, 12
                                                  30'd    4238    : data = 32'h    AFDF0B37    ;    //    lui x22 720368      ====        lui s6, 720368
                                                  30'd    4239    : data = 32'h    413DDE33    ;    //    sra x28 x27 x19      ====        sra t3, s11, s3
                                                  30'd    4240    : data = 32'h    4011D433    ;    //    sra x8 x3 x1      ====        sra s0, gp, ra
                                                  30'd    4241    : data = 32'h    0072D9B3    ;    //    srl x19 x5 x7      ====        srl s3, t0, t2
                                                  30'd    4242    : data = 32'h    00461A33    ;    //    sll x20 x12 x4      ====        sll s4, a2, tp
                                                  30'd    4243    : data = 32'h    3700CA93    ;    //    xori x21 x1 880      ====        xori s5, ra, 880
                                                  30'd    4244    : data = 32'h    0039DA13    ;    //    srli x20 x19 3      ====        srli s4, s3, 3
                                                  30'd    4245    : data = 32'h    003985B3    ;    //    add x11 x19 x3      ====        add a1, s3, gp
                                                  30'd    4246    : data = 32'h    4117DC93    ;    //    srai x25 x15 17      ====        srai s9, a5, 17
                                                  30'd    4247    : data = 32'h    007A6033    ;    //    or x0 x20 x7      ====        or zero, s4, t2
                                                  30'd    4248    : data = 32'h    E425B193    ;    //    sltiu x3 x11 -446      ====        sltiu gp, a1, -446
                                                  30'd    4249    : data = 32'h    017DE8B3    ;    //    or x17 x27 x23      ====        or a7, s11, s7
                                                  30'd    4250    : data = 32'h    01419793    ;    //    slli x15 x3 20      ====        slli a5, gp, 20
                                                  30'd    4251    : data = 32'h    0125F733    ;    //    and x14 x11 x18      ====        and a4, a1, s2
                                                  30'd    4252    : data = 32'h    34F53313    ;    //    sltiu x6 x10 847      ====        sltiu t1, a0, 847
                                                  30'd    4253    : data = 32'h    FA421B37    ;    //    lui x22 1025057      ====        lui s6, 1025057
                                                  30'd    4254    : data = 32'h    00486CB3    ;    //    or x25 x16 x4      ====        or s9, a6, tp
                                                  30'd    4255    : data = 32'h    00374D33    ;    //    xor x26 x14 x3      ====        xor s10, a4, gp
                                                  30'd    4256    : data = 32'h    CB846C13    ;    //    ori x24 x8 -840      ====        ori s8, s0, -840
                                                  30'd    4257    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4258    : data = 32'h    0DC84093    ;    //    xori x1 x16 220      ====        xori ra, a6, 220
                                                  30'd    4259    : data = 32'h    FDBA7193    ;    //    andi x3 x20 -37      ====        andi gp, s4, -37
                                                  30'd    4260    : data = 32'h    40D35B93    ;    //    srai x23 x6 13      ====        srai s7, t1, 13
                                                  30'd    4261    : data = 32'h    D2980E13    ;    //    addi x28 x16 -727      ====        addi t3, a6, -727
                                                  30'd    4262    : data = 32'h    2A9E8813    ;    //    addi x16 x29 681      ====        addi a6, t4, 681
                                                  30'd    4263    : data = 32'h    00ECA0B3    ;    //    slt x1 x25 x14      ====        slt ra, s9, a4
                                                  30'd    4264    : data = 32'h    00939D33    ;    //    sll x26 x7 x9      ====        sll s10, t2, s1
                                                  30'd    4265    : data = 32'h    017CDB33    ;    //    srl x22 x25 x23      ====        srl s6, s9, s7
                                                  30'd    4266    : data = 32'h    0012B933    ;    //    sltu x18 x5 x1      ====        sltu s2, t0, ra
                                                  30'd    4267    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4268    : data = 32'h    01AA5CB3    ;    //    srl x25 x20 x26      ====        srl s9, s4, s10
                                                  30'd    4269    : data = 32'h    00350B33    ;    //    add x22 x10 x3      ====        add s6, a0, gp
                                                  30'd    4270    : data = 32'h    32D13C13    ;    //    sltiu x24 x2 813      ====        sltiu s8, sp, 813
                                                  30'd    4271    : data = 32'h    65A7B713    ;    //    sltiu x14 x15 1626      ====        sltiu a4, a5, 1626
                                                  30'd    4272    : data = 32'h    E5992F93    ;    //    slti x31 x18 -423      ====        slti t6, s2, -423
                                                  30'd    4273    : data = 32'h    6F3F0D13    ;    //    addi x26 x30 1779      ====        addi s10, t5, 1779
                                                  30'd    4274    : data = 32'h    CFFD8293    ;    //    addi x5 x27 -769      ====        addi t0, s11, -769
                                                  30'd    4275    : data = 32'h    000E5593    ;    //    srli x11 x28 0      ====        srli a1, t3, 0
                                                  30'd    4276    : data = 32'h    62833B13    ;    //    sltiu x22 x6 1576      ====        sltiu s6, t1, 1576
                                                  30'd    4277    : data = 32'h    0071E7B3    ;    //    or x15 x3 x7      ====        or a5, gp, t2
                                                  30'd    4278    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4279    : data = 32'h    404AD1B3    ;    //    sra x3 x21 x4      ====        sra gp, s5, tp
                                                  30'd    4280    : data = 32'h    E5A50DB7    ;    //    lui x27 940624      ====        lui s11, 940624
                                                  30'd    4281    : data = 32'h    013CD5B3    ;    //    srl x11 x25 x19      ====        srl a1, s9, s3
                                                  30'd    4282    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4283    : data = 32'h    4081D9B3    ;    //    sra x19 x3 x8      ====        sra s3, gp, s0
                                                  30'd    4284    : data = 32'h    8C29B893    ;    //    sltiu x17 x19 -1854      ====        sltiu a7, s3, -1854
                                                  30'd    4285    : data = 32'h    00439393    ;    //    slli x7 x7 4      ====        slli t2, t2, 4
                                                  30'd    4286    : data = 32'h    01551D13    ;    //    slli x26 x10 21      ====        slli s10, a0, 21
                                                  30'd    4287    : data = 32'h    008735B3    ;    //    sltu x11 x14 x8      ====        sltu a1, a4, s0
                                                  30'd    4288    : data = 32'h    00E94DB3    ;    //    xor x27 x18 x14      ====        xor s11, s2, a4
                                                  30'd    4289    : data = 32'h    019945B3    ;    //    xor x11 x18 x25      ====        xor a1, s2, s9
                                                  30'd    4290    : data = 32'h    0CFF8937    ;    //    lui x18 53240      ====        lui s2, 53240
                                                  30'd    4291    : data = 32'h    00E70433    ;    //    add x8 x14 x14      ====        add s0, a4, a4
                                                  30'd    4292    : data = 32'h    4064D0B3    ;    //    sra x1 x9 x6      ====        sra ra, s1, t1
                                                  30'd    4293    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4294    : data = 32'h    7579E793    ;    //    ori x15 x19 1879      ====        ori a5, s3, 1879
                                                  30'd    4295    : data = 32'h    78196593    ;    //    ori x11 x18 1921      ====        ori a1, s2, 1921
                                                  30'd    4296    : data = 32'h    406EDD13    ;    //    srai x26 x29 6      ====        srai s10, t4, 6
                                                  30'd    4297    : data = 32'h    3F06F293    ;    //    andi x5 x13 1008      ====        andi t0, a3, 1008
                                                  30'd    4298    : data = 32'h    418ED713    ;    //    srai x14 x29 24      ====        srai a4, t4, 24
                                                  30'd    4299    : data = 32'h    01AC54B3    ;    //    srl x9 x24 x26      ====        srl s1, s8, s10
                                                  30'd    4300    : data = 32'h    06BEA293    ;    //    slti x5 x29 107      ====        slti t0, t4, 107
                                                  30'd    4301    : data = 32'h    00A67433    ;    //    and x8 x12 x10      ====        and s0, a2, a0
                                                  30'd    4302    : data = 32'h    401187B3    ;    //    sub x15 x3 x1      ====        sub a5, gp, ra
                                                  30'd    4303    : data = 32'h    9BB7D197    ;    //    auipc x3 637821      ====        auipc gp, 637821
                                                  30'd    4304    : data = 32'h    3CF36F93    ;    //    ori x31 x6 975      ====        ori t6, t1, 975
                                                  30'd    4305    : data = 32'h    09407713    ;    //    andi x14 x0 148      ====        andi a4, zero, 148
                                                  30'd    4306    : data = 32'h    7EA8A993    ;    //    slti x19 x17 2026      ====        slti s3, a7, 2026
                                                  30'd    4307    : data = 32'h    E2B48EB7    ;    //    lui x29 928584      ====        lui t4, 928584
                                                  30'd    4308    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4309    : data = 32'h    012CB8B3    ;    //    sltu x17 x25 x18      ====        sltu a7, s9, s2
                                                  30'd    4310    : data = 32'h    1AF1A037    ;    //    lui x0 110362      ====        lui zero, 110362
                                                  30'd    4311    : data = 32'h    013F5C33    ;    //    srl x24 x30 x19      ====        srl s8, t5, s3
                                                  30'd    4312    : data = 32'h    00148FB3    ;    //    add x31 x9 x1      ====        add t6, s1, ra
                                                  30'd    4313    : data = 32'h    00A2EBB3    ;    //    or x23 x5 x10      ====        or s7, t0, a0
                                                  30'd    4314    : data = 32'h    001ADEB3    ;    //    srl x29 x21 x1      ====        srl t4, s5, ra
                                                  30'd    4315    : data = 32'h    723FAC37    ;    //    lui x24 467962      ====        lui s8, 467962
                                                  30'd    4316    : data = 32'h    D013D8B7    ;    //    lui x17 852285      ====        lui a7, 852285
                                                  30'd    4317    : data = 32'h    01CBDBB3    ;    //    srl x23 x23 x28      ====        srl s7, s7, t3
                                                  30'd    4318    : data = 32'h    005F7A33    ;    //    and x20 x30 x5      ====        and s4, t5, t0
                                                  30'd    4319    : data = 32'h    F9393D13    ;    //    sltiu x26 x18 -109      ====        sltiu s10, s2, -109
                                                  30'd    4320    : data = 32'h    013ADBB3    ;    //    srl x23 x21 x19      ====        srl s7, s5, s3
                                                  30'd    4321    : data = 32'h    40248E33    ;    //    sub x28 x9 x2      ====        sub t3, s1, sp
                                                  30'd    4322    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4323    : data = 32'h    00F509B3    ;    //    add x19 x10 x15      ====        add s3, a0, a5
                                                  30'd    4324    : data = 32'h    00C7A333    ;    //    slt x6 x15 x12      ====        slt t1, a5, a2
                                                  30'd    4325    : data = 32'h    0035EFB3    ;    //    or x31 x11 x3      ====        or t6, a1, gp
                                                  30'd    4326    : data = 32'h    4E81B613    ;    //    sltiu x12 x3 1256      ====        sltiu a2, gp, 1256
                                                  30'd    4327    : data = 32'h    008EAFB3    ;    //    slt x31 x29 x8      ====        slt t6, t4, s0
                                                  30'd    4328    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4329    : data = 32'h    B787CD93    ;    //    xori x27 x15 -1160      ====        xori s11, a5, -1160
                                                  30'd    4330    : data = 32'h    00E4D433    ;    //    srl x8 x9 x14      ====        srl s0, s1, a4
                                                  30'd    4331    : data = 32'h    009B53B3    ;    //    srl x7 x22 x9      ====        srl t2, s6, s1
                                                  30'd    4332    : data = 32'h    00E45033    ;    //    srl x0 x8 x14      ====        srl zero, s0, a4
                                                  30'd    4333    : data = 32'h    6ECD8293    ;    //    addi x5 x27 1772      ====        addi t0, s11, 1772
                                                  30'd    4334    : data = 32'h    0744E013    ;    //    ori x0 x9 116      ====        ori zero, s1, 116
                                                  30'd    4335    : data = 32'h    19F82817    ;    //    auipc x16 106370      ====        auipc a6, 106370
                                                  30'd    4336    : data = 32'h    009B7FB3    ;    //    and x31 x22 x9      ====        and t6, s6, s1
                                                  30'd    4337    : data = 32'h    40BC8DB3    ;    //    sub x27 x25 x11      ====        sub s11, s9, a1
                                                  30'd    4338    : data = 32'h    0178AEB3    ;    //    slt x29 x17 x23      ====        slt t4, a7, s7
                                                  30'd    4339    : data = 32'h    01DE5E13    ;    //    srli x28 x28 29      ====        srli t3, t3, 29
                                                  30'd    4340    : data = 32'h    00DCDBB3    ;    //    srl x23 x25 x13      ====        srl s7, s9, a3
                                                  30'd    4341    : data = 32'h    7EF60713    ;    //    addi x14 x12 2031      ====        addi a4, a2, 2031
                                                  30'd    4342    : data = 32'h    017585B3    ;    //    add x11 x11 x23      ====        add a1, a1, s7
                                                  30'd    4343    : data = 32'h    1B08E593    ;    //    ori x11 x17 432      ====        ori a1, a7, 432
                                                  30'd    4344    : data = 32'h    00C8FEB3    ;    //    and x29 x17 x12      ====        and t4, a7, a2
                                                  30'd    4345    : data = 32'h    01D857B3    ;    //    srl x15 x16 x29      ====        srl a5, a6, t4
                                                  30'd    4346    : data = 32'h    43CD6413    ;    //    ori x8 x26 1084      ====        ori s0, s10, 1084
                                                  30'd    4347    : data = 32'h    2CA82813    ;    //    slti x16 x16 714      ====        slti a6, a6, 714
                                                  30'd    4348    : data = 32'h    391D2E13    ;    //    slti x28 x26 913      ====        slti t3, s10, 913
                                                  30'd    4349    : data = 32'h    01D97A33    ;    //    and x20 x18 x29      ====        and s4, s2, t4
                                                  30'd    4350    : data = 32'h    00596433    ;    //    or x8 x18 x5      ====        or s0, s2, t0
                                                  30'd    4351    : data = 32'h    40B18433    ;    //    sub x8 x3 x11      ====        sub s0, gp, a1
                                                  30'd    4352    : data = 32'h    01CD91B3    ;    //    sll x3 x27 x28      ====        sll gp, s11, t3
                                                  30'd    4353    : data = 32'h    0D0D7193    ;    //    andi x3 x26 208      ====        andi gp, s10, 208
                                                  30'd    4354    : data = 32'h    00427033    ;    //    and x0 x4 x4      ====        and zero, tp, tp
                                                  30'd    4355    : data = 32'h    5F438A97    ;    //    auipc x21 390200      ====        auipc s5, 390200
                                                  30'd    4356    : data = 32'h    E63D5B97    ;    //    auipc x23 943061      ====        auipc s7, 943061
                                                  30'd    4357    : data = 32'h    D565F137    ;    //    lui x2 874079      ====        lui sp, 874079
                                                  30'd    4358    : data = 32'h    71DF4A93    ;    //    xori x21 x30 1821      ====        xori s5, t5, 1821
                                                  30'd    4359    : data = 32'h    005582B3    ;    //    add x5 x11 x5      ====        add t0, a1, t0
                                                  30'd    4360    : data = 32'h    01FDD0B3    ;    //    srl x1 x27 x31      ====        srl ra, s11, t6
                                                  30'd    4361    : data = 32'h    665F4497    ;    //    auipc x9 419316      ====        auipc s1, 419316
                                                  30'd    4362    : data = 32'h    40BED013    ;    //    srai x0 x29 11      ====        srai zero, t4, 11
                                                  30'd    4363    : data = 32'h    0967E993    ;    //    ori x19 x15 150      ====        ori s3, a5, 150
                                                  30'd    4364    : data = 32'h    9B628117    ;    //    auipc x2 636456      ====        auipc sp, 636456
                                                  30'd    4365    : data = 32'h    970DF5B7    ;    //    lui x11 618719      ====        lui a1, 618719
                                                  30'd    4366    : data = 32'h    A012CD17    ;    //    auipc x26 655660      ====        auipc s10, 655660
                                                  30'd    4367    : data = 32'h    C6166993    ;    //    ori x19 x12 -927      ====        ori s3, a2, -927
                                                  30'd    4368    : data = 32'h    C2162293    ;    //    slti x5 x12 -991      ====        slti t0, a2, -991
                                                  30'd    4369    : data = 32'h    5D8E6713    ;    //    ori x14 x28 1496      ====        ori a4, t3, 1496
                                                  30'd    4370    : data = 32'h    007B9793    ;    //    slli x15 x23 7      ====        slli a5, s7, 7
                                                  30'd    4371    : data = 32'h    41F68AB3    ;    //    sub x21 x13 x31      ====        sub s5, a3, t6
                                                  30'd    4372    : data = 32'h    010DE4B3    ;    //    or x9 x27 x16      ====        or s1, s11, a6
                                                  30'd    4373    : data = 32'h    0E2A6013    ;    //    ori x0 x20 226      ====        ori zero, s4, 226
                                                  30'd    4374    : data = 32'h    0115BFB3    ;    //    sltu x31 x11 x17      ====        sltu t6, a1, a7
                                                  30'd    4375    : data = 32'h    4092DD93    ;    //    srai x27 x5 9      ====        srai s11, t0, 9
                                                  30'd    4376    : data = 32'h    00CCF133    ;    //    and x2 x25 x12      ====        and sp, s9, a2
                                                  30'd    4377    : data = 32'h    01A61333    ;    //    sll x6 x12 x26      ====        sll t1, a2, s10
                                                  30'd    4378    : data = 32'h    98CCEC13    ;    //    ori x24 x25 -1652      ====        ori s8, s9, -1652
                                                  30'd    4379    : data = 32'h    95CC7113    ;    //    andi x2 x24 -1700      ====        andi sp, s8, -1700
                                                  30'd    4380    : data = 32'h    4048D833    ;    //    sra x16 x17 x4      ====        sra a6, a7, tp
                                                  30'd    4381    : data = 32'h    DFB17E13    ;    //    andi x28 x2 -517      ====        andi t3, sp, -517
                                                  30'd    4382    : data = 32'h    00BA34B3    ;    //    sltu x9 x20 x11      ====        sltu s1, s4, a1
                                                  30'd    4383    : data = 32'h    010AF8B3    ;    //    and x17 x21 x16      ====        and a7, s5, a6
                                                  30'd    4384    : data = 32'h    E1FF3613    ;    //    sltiu x12 x30 -481      ====        sltiu a2, t5, -481
                                                  30'd    4385    : data = 32'h    7A1C0497    ;    //    auipc x9 500160      ====        auipc s1, 500160
                                                  30'd    4386    : data = 32'h    01716E33    ;    //    or x28 x2 x23      ====        or t3, sp, s7
                                                  30'd    4387    : data = 32'h    00D3DCB3    ;    //    srl x25 x7 x13      ====        srl s9, t2, a3
                                                  30'd    4388    : data = 32'h    3E74A637    ;    //    lui x12 255818      ====        lui a2, 255818
                                                  30'd    4389    : data = 32'h    F6333613    ;    //    sltiu x12 x6 -157      ====        sltiu a2, t1, -157
                                                  30'd    4390    : data = 32'h    01845393    ;    //    srli x7 x8 24      ====        srli t2, s0, 24
                                                  30'd    4391    : data = 32'h    AA111697    ;    //    auipc x13 696593      ====        auipc a3, 696593
                                                  30'd    4392    : data = 32'h    B3A7C313    ;    //    xori x6 x15 -1222      ====        xori t1, a5, -1222
                                                  30'd    4393    : data = 32'h    0114D3B3    ;    //    srl x7 x9 x17      ====        srl t2, s1, a7
                                                  30'd    4394    : data = 32'h    40EFDAB3    ;    //    sra x21 x31 x14      ====        sra s5, t6, a4
                                                  30'd    4395    : data = 32'h    D361DF97    ;    //    auipc x31 865821      ====        auipc t6, 865821
                                                  30'd    4396    : data = 32'h    01A71AB3    ;    //    sll x21 x14 x26      ====        sll s5, a4, s10
                                                  30'd    4397    : data = 32'h    733AF813    ;    //    andi x16 x21 1843      ====        andi a6, s5, 1843
                                                  30'd    4398    : data = 32'h    0C22CA93    ;    //    xori x21 x5 194      ====        xori s5, t0, 194
                                                  30'd    4399    : data = 32'h    006FD613    ;    //    srli x12 x31 6      ====        srli a2, t6, 6
                                                  30'd    4400    : data = 32'h    017482B3    ;    //    add x5 x9 x23      ====        add t0, s1, s7
                                                  30'd    4401    : data = 32'h    00B23833    ;    //    sltu x16 x4 x11      ====        sltu a6, tp, a1
                                                  30'd    4402    : data = 32'h    671F0993    ;    //    addi x19 x30 1649      ====        addi s3, t5, 1649
                                                  30'd    4403    : data = 32'h    014532B3    ;    //    sltu x5 x10 x20      ====        sltu t0, a0, s4
                                                  30'd    4404    : data = 32'h    01068133    ;    //    add x2 x13 x16      ====        add sp, a3, a6
                                                  30'd    4405    : data = 32'h    AFB33713    ;    //    sltiu x14 x6 -1285      ====        sltiu a4, t1, -1285
                                                  30'd    4406    : data = 32'h    406DD333    ;    //    sra x6 x27 x6      ====        sra t1, s11, t1
                                                  30'd    4407    : data = 32'h    0060BA33    ;    //    sltu x20 x1 x6      ====        sltu s4, ra, t1
                                                  30'd    4408    : data = 32'h    1DE74693    ;    //    xori x13 x14 478      ====        xori a3, a4, 478
                                                  30'd    4409    : data = 32'h    00A2BDB3    ;    //    sltu x27 x5 x10      ====        sltu s11, t0, a0
                                                  30'd    4410    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4411    : data = 32'h    17200193    ;    //    addi x3 x0 370      ====        addi gp, zero, 370
                                                  30'd    4412    : data = 32'h    007FDFB3    ;    //    srl x31 x31 x7      ====        srl t6, t6, t2
                                                  30'd    4413    : data = 32'h    E99F7993    ;    //    andi x19 x30 -359      ====        andi s3, t5, -359
                                                  30'd    4414    : data = 32'h    41D08633    ;    //    sub x12 x1 x29      ====        sub a2, ra, t4
                                                  30'd    4415    : data = 32'h    00551713    ;    //    slli x14 x10 5      ====        slli a4, a0, 5
                                                  30'd    4416    : data = 32'h    4141D013    ;    //    srai x0 x3 20      ====        srai zero, gp, 20
                                                  30'd    4417    : data = 32'h    01FB7B33    ;    //    and x22 x22 x31      ====        and s6, s6, t6
                                                  30'd    4418    : data = 32'h    498B2C93    ;    //    slti x25 x22 1176      ====        slti s9, s6, 1176
                                                  30'd    4419    : data = 32'h    016D0433    ;    //    add x8 x26 x22      ====        add s0, s10, s6
                                                  30'd    4420    : data = 32'h    41315D13    ;    //    srai x26 x2 19      ====        srai s10, sp, 19
                                                  30'd    4421    : data = 32'h    7FCDE113    ;    //    ori x2 x27 2044      ====        ori sp, s11, 2044
                                                  30'd    4422    : data = 32'h    00F1BD33    ;    //    sltu x26 x3 x15      ====        sltu s10, gp, a5
                                                  30'd    4423    : data = 32'h    00678EB3    ;    //    add x29 x15 x6      ====        add t4, a5, t1
                                                  30'd    4424    : data = 32'h    009D2D33    ;    //    slt x26 x26 x9      ====        slt s10, s10, s1
                                                  30'd    4425    : data = 32'h    017C5193    ;    //    srli x3 x24 23      ====        srli gp, s8, 23
                                                  30'd    4426    : data = 32'h    F67D8A13    ;    //    addi x20 x27 -153      ====        addi s4, s11, -153
                                                  30'd    4427    : data = 32'h    F5BCC2B7    ;    //    lui x5 1006540      ====        lui t0, 1006540
                                                  30'd    4428    : data = 32'h    00E6ECB3    ;    //    or x25 x13 x14      ====        or s9, a3, a4
                                                  30'd    4429    : data = 32'h    E96E6113    ;    //    ori x2 x28 -362      ====        ori sp, t3, -362
                                                  30'd    4430    : data = 32'h    95AB7D93    ;    //    andi x27 x22 -1702      ====        andi s11, s6, -1702
                                                  30'd    4431    : data = 32'h    017969B3    ;    //    or x19 x18 x23      ====        or s3, s2, s7
                                                  30'd    4432    : data = 32'h    00A6E1B3    ;    //    or x3 x13 x10      ====        or gp, a3, a0
                                                  30'd    4433    : data = 32'h    01277033    ;    //    and x0 x14 x18      ====        and zero, a4, s2
                                                  30'd    4434    : data = 32'h    A4F09437    ;    //    lui x8 675593      ====        lui s0, 675593
                                                  30'd    4435    : data = 32'h    41A583B3    ;    //    sub x7 x11 x26      ====        sub t2, a1, s10
                                                  30'd    4436    : data = 32'h    41BBDF93    ;    //    srai x31 x23 27      ====        srai t6, s7, 27
                                                  30'd    4437    : data = 32'h    6235AC13    ;    //    slti x24 x11 1571      ====        slti s8, a1, 1571
                                                  30'd    4438    : data = 32'h    0199E7B3    ;    //    or x15 x19 x25      ====        or a5, s3, s9
                                                  30'd    4439    : data = 32'h    00CC3833    ;    //    sltu x16 x24 x12      ====        sltu a6, s8, a2
                                                  30'd    4440    : data = 32'h    0194D093    ;    //    srli x1 x9 25      ====        srli ra, s1, 25
                                                  30'd    4441    : data = 32'h    00854E33    ;    //    xor x28 x10 x8      ====        xor t3, a0, s0
                                                  30'd    4442    : data = 32'h    004E18B3    ;    //    sll x17 x28 x4      ====        sll a7, t3, tp
                                                  30'd    4443    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4444    : data = 32'h    AE7AE493    ;    //    ori x9 x21 -1305      ====        ori s1, s5, -1305
                                                  30'd    4445    : data = 32'h    55357993    ;    //    andi x19 x10 1363      ====        andi s3, a0, 1363
                                                  30'd    4446    : data = 32'h    01E64DB3    ;    //    xor x27 x12 x30      ====        xor s11, a2, t5
                                                  30'd    4447    : data = 32'h    40E303B3    ;    //    sub x7 x6 x14      ====        sub t2, t1, a4
                                                  30'd    4448    : data = 32'h    00277833    ;    //    and x16 x14 x2      ====        and a6, a4, sp
                                                  30'd    4449    : data = 32'h    5ACE6293    ;    //    ori x5 x28 1452      ====        ori t0, t3, 1452
                                                  30'd    4450    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4451    : data = 32'h    018DF9B3    ;    //    and x19 x27 x24      ====        and s3, s11, s8
                                                  30'd    4452    : data = 32'h    00474BB3    ;    //    xor x23 x14 x4      ====        xor s7, a4, tp
                                                  30'd    4453    : data = 32'h    0007D6B3    ;    //    srl x13 x15 x0      ====        srl a3, a5, zero
                                                  30'd    4454    : data = 32'h    01DB9A33    ;    //    sll x20 x23 x29      ====        sll s4, s7, t4
                                                  30'd    4455    : data = 32'h    01A25813    ;    //    srli x16 x4 26      ====        srli a6, tp, 26
                                                  30'd    4456    : data = 32'h    00DA0833    ;    //    add x16 x20 x13      ====        add a6, s4, a3
                                                  30'd    4457    : data = 32'h    BABA7293    ;    //    andi x5 x20 -1109      ====        andi t0, s4, -1109
                                                  30'd    4458    : data = 32'h    0128CCB3    ;    //    xor x25 x17 x18      ====        xor s9, a7, s2
                                                  30'd    4459    : data = 32'h    011E5393    ;    //    srli x7 x28 17      ====        srli t2, t3, 17
                                                  30'd    4460    : data = 32'h    416C5313    ;    //    srai x6 x24 22      ====        srai t1, s8, 22
                                                  30'd    4461    : data = 32'h    00589733    ;    //    sll x14 x17 x5      ====        sll a4, a7, t0
                                                  30'd    4462    : data = 32'h    31132D13    ;    //    slti x26 x6 785      ====        slti s10, t1, 785
                                                  30'd    4463    : data = 32'h    0031E133    ;    //    or x2 x3 x3      ====        or sp, gp, gp
                                                  30'd    4464    : data = 32'h    00409913    ;    //    slli x18 x1 4      ====        slli s2, ra, 4
                                                  30'd    4465    : data = 32'h    01448433    ;    //    add x8 x9 x20      ====        add s0, s1, s4
                                                  30'd    4466    : data = 32'h    0098F8B3    ;    //    and x17 x17 x9      ====        and a7, a7, s1
                                                  30'd    4467    : data = 32'h    413E5713    ;    //    srai x14 x28 19      ====        srai a4, t3, 19
                                                  30'd    4468    : data = 32'h    005D5E33    ;    //    srl x28 x26 x5      ====        srl t3, s10, t0
                                                  30'd    4469    : data = 32'h    40CE7393    ;    //    andi x7 x28 1036      ====        andi t2, t3, 1036
                                                  30'd    4470    : data = 32'h    01495393    ;    //    srli x7 x18 20      ====        srli t2, s2, 20
                                                  30'd    4471    : data = 32'h    9E086993    ;    //    ori x19 x16 -1568      ====        ori s3, a6, -1568
                                                  30'd    4472    : data = 32'h    0109B1B3    ;    //    sltu x3 x19 x16      ====        sltu gp, s3, a6
                                                  30'd    4473    : data = 32'h    40A35493    ;    //    srai x9 x6 10      ====        srai s1, t1, 10
                                                  30'd    4474    : data = 32'h    FCD9CB93    ;    //    xori x23 x19 -51      ====        xori s7, s3, -51
                                                  30'd    4475    : data = 32'h    01678833    ;    //    add x16 x15 x22      ====        add a6, a5, s6
                                                  30'd    4476    : data = 32'h    D6BE7EB7    ;    //    lui x29 879591      ====        lui t4, 879591
                                                  30'd    4477    : data = 32'h    01D782B3    ;    //    add x5 x15 x29      ====        add t0, a5, t4
                                                  30'd    4478    : data = 32'h    01241493    ;    //    slli x9 x8 18      ====        slli s1, s0, 18
                                                  30'd    4479    : data = 32'h    C998EB93    ;    //    ori x23 x17 -871      ====        ori s7, a7, -871
                                                  30'd    4480    : data = 32'h    40ACDD13    ;    //    srai x26 x25 10      ====        srai s10, s9, 10
                                                  30'd    4481    : data = 32'h    BC2C4993    ;    //    xori x19 x24 -1086      ====        xori s3, s8, -1086
                                                  30'd    4482    : data = 32'h    00AFD693    ;    //    srli x13 x31 10      ====        srli a3, t6, 10
                                                  30'd    4483    : data = 32'h    41D006B3    ;    //    sub x13 x0 x29      ====        sub a3, zero, t4
                                                  30'd    4484    : data = 32'h    40000FB3    ;    //    sub x31 x0 x0      ====        sub t6, zero, zero
                                                  30'd    4485    : data = 32'h    00786733    ;    //    or x14 x16 x7      ====        or a4, a6, t2
                                                  30'd    4486    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4487    : data = 32'h    0DD21137    ;    //    lui x2 56609      ====        lui sp, 56609
                                                  30'd    4488    : data = 32'h    A548B113    ;    //    sltiu x2 x17 -1452      ====        sltiu sp, a7, -1452
                                                  30'd    4489    : data = 32'h    957A8893    ;    //    addi x17 x21 -1705      ====        addi a7, s5, -1705
                                                  30'd    4490    : data = 32'h    162BB593    ;    //    sltiu x11 x23 354      ====        sltiu a1, s7, 354
                                                  30'd    4491    : data = 32'h    0094DC33    ;    //    srl x24 x9 x9      ====        srl s8, s1, s1
                                                  30'd    4492    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4493    : data = 32'h    410A0633    ;    //    sub x12 x20 x16      ====        sub a2, s4, a6
                                                  30'd    4494    : data = 32'h    00B6ABB3    ;    //    slt x23 x13 x11      ====        slt s7, a3, a1
                                                  30'd    4495    : data = 32'h    4031D133    ;    //    sra x2 x3 x3      ====        sra sp, gp, gp
                                                  30'd    4496    : data = 32'h    00AE1E13    ;    //    slli x28 x28 10      ====        slli t3, t3, 10
                                                  30'd    4497    : data = 32'h    182BC713    ;    //    xori x14 x23 386      ====        xori a4, s7, 386
                                                  30'd    4498    : data = 32'h    01F53FB3    ;    //    sltu x31 x10 x31      ====        sltu t6, a0, t6
                                                  30'd    4499    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4500    : data = 32'h    F2316593    ;    //    ori x11 x2 -221      ====        ori a1, sp, -221
                                                  30'd    4501    : data = 32'h    002537B3    ;    //    sltu x15 x10 x2      ====        sltu a5, a0, sp
                                                  30'd    4502    : data = 32'h    00681F93    ;    //    slli x31 x16 6      ====        slli t6, a6, 6
                                                  30'd    4503    : data = 32'h    01BE22B3    ;    //    slt x5 x28 x27      ====        slt t0, t3, s11
                                                  30'd    4504    : data = 32'h    1D2D3C13    ;    //    sltiu x24 x26 466      ====        sltiu s8, s10, 466
                                                  30'd    4505    : data = 32'h    01F0EA33    ;    //    or x20 x1 x31      ====        or s4, ra, t6
                                                  30'd    4506    : data = 32'h    41C58D33    ;    //    sub x26 x11 x28      ====        sub s10, a1, t3
                                                  30'd    4507    : data = 32'h    462EA6B7    ;    //    lui x13 287466      ====        lui a3, 287466
                                                  30'd    4508    : data = 32'h    40CEDC93    ;    //    srai x25 x29 12      ====        srai s9, t4, 12
                                                  30'd    4509    : data = 32'h    D59D3793    ;    //    sltiu x15 x26 -679      ====        sltiu a5, s10, -679
                                                  30'd    4510    : data = 32'h    41A3DA33    ;    //    sra x20 x7 x26      ====        sra s4, t2, s10
                                                  30'd    4511    : data = 32'h    00E325B3    ;    //    slt x11 x6 x14      ====        slt a1, t1, a4
                                                  30'd    4512    : data = 32'h    A9F2F193    ;    //    andi x3 x5 -1377      ====        andi gp, t0, -1377
                                                  30'd    4513    : data = 32'h    01214033    ;    //    xor x0 x2 x18      ====        xor zero, sp, s2
                                                  30'd    4514    : data = 32'h    00BA7033    ;    //    and x0 x20 x11      ====        and zero, s4, a1
                                                  30'd    4515    : data = 32'h    00AD2FB3    ;    //    slt x31 x26 x10      ====        slt t6, s10, a0
                                                  30'd    4516    : data = 32'h    00D580B3    ;    //    add x1 x11 x13      ====        add ra, a1, a3
                                                  30'd    4517    : data = 32'h    568A3D13    ;    //    sltiu x26 x20 1384      ====        sltiu s10, s4, 1384
                                                  30'd    4518    : data = 32'h    40D2D033    ;    //    sra x0 x5 x13      ====        sra zero, t0, a3
                                                  30'd    4519    : data = 32'h    01314DB3    ;    //    xor x27 x2 x19      ====        xor s11, sp, s3
                                                  30'd    4520    : data = 32'h    00831993    ;    //    slli x19 x6 8      ====        slli s3, t1, 8
                                                  30'd    4521    : data = 32'h    7D0F3117    ;    //    auipc x2 512243      ====        auipc sp, 512243
                                                  30'd    4522    : data = 32'h    01AC23B3    ;    //    slt x7 x24 x26      ====        slt t2, s8, s10
                                                  30'd    4523    : data = 32'h    009C15B3    ;    //    sll x11 x24 x9      ====        sll a1, s8, s1
                                                  30'd    4524    : data = 32'h    00791293    ;    //    slli x5 x18 7      ====        slli t0, s2, 7
                                                  30'd    4525    : data = 32'h    18036293    ;    //    ori x5 x6 384      ====        ori t0, t1, 384
                                                  30'd    4526    : data = 32'h    01648E33    ;    //    add x28 x9 x22      ====        add t3, s1, s6
                                                  30'd    4527    : data = 32'h    8CD66813    ;    //    ori x16 x12 -1843      ====        ori a6, a2, -1843
                                                  30'd    4528    : data = 32'h    EA9E4013    ;    //    xori x0 x28 -343      ====        xori zero, t3, -343
                                                  30'd    4529    : data = 32'h    01CDDC93    ;    //    srli x25 x27 28      ====        srli s9, s11, 28
                                                  30'd    4530    : data = 32'h    01147B33    ;    //    and x22 x8 x17      ====        and s6, s0, a7
                                                  30'd    4531    : data = 32'h    F126CE93    ;    //    xori x29 x13 -238      ====        xori t4, a3, -238
                                                  30'd    4532    : data = 32'h    01C32033    ;    //    slt x0 x6 x28      ====        slt zero, t1, t3
                                                  30'd    4533    : data = 32'h    6B013D13    ;    //    sltiu x26 x2 1712      ====        sltiu s10, sp, 1712
                                                  30'd    4534    : data = 32'h    83764413    ;    //    xori x8 x12 -1993      ====        xori s0, a2, -1993
                                                  30'd    4535    : data = 32'h    2C66C813    ;    //    xori x16 x13 710      ====        xori a6, a3, 710
                                                  30'd    4536    : data = 32'h    4117D913    ;    //    srai x18 x15 17      ====        srai s2, a5, 17
                                                  30'd    4537    : data = 32'h    C54AA393    ;    //    slti x7 x21 -940      ====        slti t2, s5, -940
                                                  30'd    4538    : data = 32'h    00117FB3    ;    //    and x31 x2 x1      ====        and t6, sp, ra
                                                  30'd    4539    : data = 32'h    401DD9B3    ;    //    sra x19 x27 x1      ====        sra s3, s11, ra
                                                  30'd    4540    : data = 32'h    01CB5113    ;    //    srli x2 x22 28      ====        srli sp, s6, 28
                                                  30'd    4541    : data = 32'h    00ADEDB3    ;    //    or x27 x27 x10      ====        or s11, s11, a0
                                                  30'd    4542    : data = 32'h    0069B833    ;    //    sltu x16 x19 x6      ====        sltu a6, s3, t1
                                                  30'd    4543    : data = 32'h    0048D713    ;    //    srli x14 x17 4      ====        srli a4, a7, 4
                                                  30'd    4544    : data = 32'h    B4C5BDB7    ;    //    lui x27 740443      ====        lui s11, 740443
                                                  30'd    4545    : data = 32'h    41CCDCB3    ;    //    sra x25 x25 x28      ====        sra s9, s9, t3
                                                  30'd    4546    : data = 32'h    3D9F3A93    ;    //    sltiu x21 x30 985      ====        sltiu s5, t5, 985
                                                  30'd    4547    : data = 32'h    0029BE33    ;    //    sltu x28 x19 x2      ====        sltu t3, s3, sp
                                                  30'd    4548    : data = 32'h    01375A93    ;    //    srli x21 x14 19      ====        srli s5, a4, 19
                                                  30'd    4549    : data = 32'h    01847733    ;    //    and x14 x8 x24      ====        and a4, s0, s8
                                                  30'd    4550    : data = 32'h    FC75FD13    ;    //    andi x26 x11 -57      ====        andi s10, a1, -57
                                                  30'd    4551    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4552    : data = 32'h    188C4E17    ;    //    auipc x28 100548      ====        auipc t3, 100548
                                                  30'd    4553    : data = 32'h    FA438A93    ;    //    addi x21 x7 -92      ====        addi s5, t2, -92
                                                  30'd    4554    : data = 32'h    36DA8193    ;    //    addi x3 x21 877      ====        addi gp, s5, 877
                                                  30'd    4555    : data = 32'h    008C1FB3    ;    //    sll x31 x24 x8      ====        sll t6, s8, s0
                                                  30'd    4556    : data = 32'h    DDF1BD13    ;    //    sltiu x26 x3 -545      ====        sltiu s10, gp, -545
                                                  30'd    4557    : data = 32'h    8D0ECC13    ;    //    xori x24 x29 -1840      ====        xori s8, t4, -1840
                                                  30'd    4558    : data = 32'h    010283B3    ;    //    add x7 x5 x16      ====        add t2, t0, a6
                                                  30'd    4559    : data = 32'h    74D67D37    ;    //    lui x26 478567      ====        lui s10, 478567
                                                  30'd    4560    : data = 32'h    01551693    ;    //    slli x13 x10 21      ====        slli a3, a0, 21
                                                  30'd    4561    : data = 32'h    01DCD093    ;    //    srli x1 x25 29      ====        srli ra, s9, 29
                                                  30'd    4562    : data = 32'h    411FDC13    ;    //    srai x24 x31 17      ====        srai s8, t6, 17
                                                  30'd    4563    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4564    : data = 32'h    405CD193    ;    //    srai x3 x25 5      ====        srai gp, s9, 5
                                                  30'd    4565    : data = 32'h    01BB3033    ;    //    sltu x0 x22 x27      ====        sltu zero, s6, s11
                                                  30'd    4566    : data = 32'h    DEF3AA13    ;    //    slti x20 x7 -529      ====        slti s4, t2, -529
                                                  30'd    4567    : data = 32'h    673B2393    ;    //    slti x7 x22 1651      ====        slti t2, s6, 1651
                                                  30'd    4568    : data = 32'h    001FF733    ;    //    and x14 x31 x1      ====        and a4, t6, ra
                                                  30'd    4569    : data = 32'h    279C0E13    ;    //    addi x28 x24 633      ====        addi t3, s8, 633
                                                  30'd    4570    : data = 32'h    01451C93    ;    //    slli x25 x10 20      ====        slli s9, a0, 20
                                                  30'd    4571    : data = 32'h    00F01EB3    ;    //    sll x29 x0 x15      ====        sll t4, zero, a5
                                                  30'd    4572    : data = 32'h    40FF5A13    ;    //    srai x20 x30 15      ====        srai s4, t5, 15
                                                  30'd    4573    : data = 32'h    2DAB3493    ;    //    sltiu x9 x22 730      ====        sltiu s1, s6, 730
                                                  30'd    4574    : data = 32'h    41B305B3    ;    //    sub x11 x6 x27      ====        sub a1, t1, s11
                                                  30'd    4575    : data = 32'h    01B7E833    ;    //    or x16 x15 x27      ====        or a6, a5, s11
                                                  30'd    4576    : data = 32'h    00F89833    ;    //    sll x16 x17 x15      ====        sll a6, a7, a5
                                                  30'd    4577    : data = 32'h    12467D13    ;    //    andi x26 x12 292      ====        andi s10, a2, 292
                                                  30'd    4578    : data = 32'h    00BD80B3    ;    //    add x1 x27 x11      ====        add ra, s11, a1
                                                  30'd    4579    : data = 32'h    829CB893    ;    //    sltiu x17 x25 -2007      ====        sltiu a7, s9, -2007
                                                  30'd    4580    : data = 32'h    01900D33    ;    //    add x26 x0 x25      ====        add s10, zero, s9
                                                  30'd    4581    : data = 32'h    002FB1B3    ;    //    sltu x3 x31 x2      ====        sltu gp, t6, sp
                                                  30'd    4582    : data = 32'h    01AF9133    ;    //    sll x2 x31 x26      ====        sll sp, t6, s10
                                                  30'd    4583    : data = 32'h    CBF9C713    ;    //    xori x14 x19 -833      ====        xori a4, s3, -833
                                                  30'd    4584    : data = 32'h    00AA5B13    ;    //    srli x22 x20 10      ====        srli s6, s4, 10
                                                  30'd    4585    : data = 32'h    014ED8B3    ;    //    srl x17 x29 x20      ====        srl a7, t4, s4
                                                  30'd    4586    : data = 32'h    01C25193    ;    //    srli x3 x4 28      ====        srli gp, tp, 28
                                                  30'd    4587    : data = 32'h    7C763E37    ;    //    lui x28 509795      ====        lui t3, 509795
                                                  30'd    4588    : data = 32'h    B4757D17    ;    //    auipc x26 739159      ====        auipc s10, 739159
                                                  30'd    4589    : data = 32'h    E07F8993    ;    //    addi x19 x31 -505      ====        addi s3, t6, -505
                                                  30'd    4590    : data = 32'h    CA34BC13    ;    //    sltiu x24 x9 -861      ====        sltiu s8, s1, -861
                                                  30'd    4591    : data = 32'h    00CBF0B3    ;    //    and x1 x23 x12      ====        and ra, s7, a2
                                                  30'd    4592    : data = 32'h    A66C2193    ;    //    slti x3 x24 -1434      ====        slti gp, s8, -1434
                                                  30'd    4593    : data = 32'h    00DB3C33    ;    //    sltu x24 x22 x13      ====        sltu s8, s6, a3
                                                  30'd    4594    : data = 32'h    E9C4AB13    ;    //    slti x22 x9 -356      ====        slti s6, s1, -356
                                                  30'd    4595    : data = 32'h    4064D713    ;    //    srai x14 x9 6      ====        srai a4, s1, 6
                                                  30'd    4596    : data = 32'h    05382013    ;    //    slti x0 x16 83      ====        slti zero, a6, 83
                                                  30'd    4597    : data = 32'h    8C200B93    ;    //    addi x23 x0 -1854      ====        addi s7, zero, -1854
                                                  30'd    4598    : data = 32'h    01FDD733    ;    //    srl x14 x27 x31      ====        srl a4, s11, t6
                                                  30'd    4599    : data = 32'h    F9B86E13    ;    //    ori x28 x16 -101      ====        ori t3, a6, -101
                                                  30'd    4600    : data = 32'h    CF73AD93    ;    //    slti x27 x7 -777      ====        slti s11, t2, -777
                                                  30'd    4601    : data = 32'h    4152DD93    ;    //    srai x27 x5 21      ====        srai s11, t0, 21
                                                  30'd    4602    : data = 32'h    01603D33    ;    //    sltu x26 x0 x22      ====        sltu s10, zero, s6
                                                  30'd    4603    : data = 32'h    BE1A2913    ;    //    slti x18 x20 -1055      ====        slti s2, s4, -1055
                                                  30'd    4604    : data = 32'h    F20FC997    ;    //    auipc x19 991484      ====        auipc s3, 991484
                                                  30'd    4605    : data = 32'h    01401493    ;    //    slli x9 x0 20      ====        slli s1, zero, 20
                                                  30'd    4606    : data = 32'h    00624033    ;    //    xor x0 x4 x6      ====        xor zero, tp, t1
                                                  30'd    4607    : data = 32'h    21F82D93    ;    //    slti x27 x16 543      ====        slti s11, a6, 543
                                                  30'd    4608    : data = 32'h    4353F313    ;    //    andi x6 x7 1077      ====        andi t1, t2, 1077
                                                  30'd    4609    : data = 32'h    0131EC33    ;    //    or x24 x3 x19      ====        or s8, gp, s3
                                                  30'd    4610    : data = 32'h    01880133    ;    //    add x2 x16 x24      ====        add sp, a6, s8
                                                  30'd    4611    : data = 32'h    013B12B3    ;    //    sll x5 x22 x19      ====        sll t0, s6, s3
                                                  30'd    4612    : data = 32'h    000D5333    ;    //    srl x6 x26 x0      ====        srl t1, s10, zero
                                                  30'd    4613    : data = 32'h    07074713    ;    //    xori x14 x14 112      ====        xori a4, a4, 112
                                                  30'd    4614    : data = 32'h    40420A33    ;    //    sub x20 x4 x4      ====        sub s4, tp, tp
                                                  30'd    4615    : data = 32'h    9CC59737    ;    //    lui x14 642137      ====        lui a4, 642137
                                                  30'd    4616    : data = 32'h    B1270397    ;    //    auipc x7 725616      ====        auipc t2, 725616
                                                  30'd    4617    : data = 32'h    000B5493    ;    //    srli x9 x22 0      ====        srli s1, s6, 0
                                                  30'd    4618    : data = 32'h    2ECB2617    ;    //    auipc x12 191666      ====        auipc a2, 191666
                                                  30'd    4619    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4620    : data = 32'h    0003FBB3    ;    //    and x23 x7 x0      ====        and s7, t2, zero
                                                  30'd    4621    : data = 32'h    0180DB93    ;    //    srli x23 x1 24      ====        srli s7, ra, 24
                                                  30'd    4622    : data = 32'h    40C55433    ;    //    sra x8 x10 x12      ====        sra s0, a0, a2
                                                  30'd    4623    : data = 32'h    002BFFB3    ;    //    and x31 x23 x2      ====        and t6, s7, sp
                                                  30'd    4624    : data = 32'h    001E25B3    ;    //    slt x11 x28 x1      ====        slt a1, t3, ra
                                                  30'd    4625    : data = 32'h    D0257437    ;    //    lui x8 852567      ====        lui s0, 852567
                                                  30'd    4626    : data = 32'h    577DE713    ;    //    ori x14 x27 1399      ====        ori a4, s11, 1399
                                                  30'd    4627    : data = 32'h    40B2DB33    ;    //    sra x22 x5 x11      ====        sra s6, t0, a1
                                                  30'd    4628    : data = 32'h    01BD5B33    ;    //    srl x22 x26 x27      ====        srl s6, s10, s11
                                                  30'd    4629    : data = 32'h    B76FF613    ;    //    andi x12 x31 -1162      ====        andi a2, t6, -1162
                                                  30'd    4630    : data = 32'h    016E1C33    ;    //    sll x24 x28 x22      ====        sll s8, t3, s6
                                                  30'd    4631    : data = 32'h    01DA85B3    ;    //    add x11 x21 x29      ====        add a1, s5, t4
                                                  30'd    4632    : data = 32'h    003130B3    ;    //    sltu x1 x2 x3      ====        sltu ra, sp, gp
                                                  30'd    4633    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4634    : data = 32'h    016926B3    ;    //    slt x13 x18 x22      ====        slt a3, s2, s6
                                                  30'd    4635    : data = 32'h    004C2D33    ;    //    slt x26 x24 x4      ====        slt s10, s8, tp
                                                  30'd    4636    : data = 32'h    01557133    ;    //    and x2 x10 x21      ====        and sp, a0, s5
                                                  30'd    4637    : data = 32'h    459DBE93    ;    //    sltiu x29 x27 1113      ====        sltiu t4, s11, 1113
                                                  30'd    4638    : data = 32'h    00CC54B3    ;    //    srl x9 x24 x12      ====        srl s1, s8, a2
                                                  30'd    4639    : data = 32'h    D8464E37    ;    //    lui x28 885860      ====        lui t3, 885860
                                                  30'd    4640    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4641    : data = 32'h    D9188013    ;    //    addi x0 x17 -623      ====        addi zero, a7, -623
                                                  30'd    4642    : data = 32'h    C0382B13    ;    //    slti x22 x16 -1021      ====        slti s6, a6, -1021
                                                  30'd    4643    : data = 32'h    04A72393    ;    //    slti x7 x14 74      ====        slti t2, a4, 74
                                                  30'd    4644    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4645    : data = 32'h    40485593    ;    //    srai x11 x16 4      ====        srai a1, a6, 4
                                                  30'd    4646    : data = 32'h    01B303B3    ;    //    add x7 x6 x27      ====        add t2, t1, s11
                                                  30'd    4647    : data = 32'h    0087F3B3    ;    //    and x7 x15 x8      ====        and t2, a5, s0
                                                  30'd    4648    : data = 32'h    00DC3A33    ;    //    sltu x20 x24 x13      ====        sltu s4, s8, a3
                                                  30'd    4649    : data = 32'h    4019D313    ;    //    srai x6 x19 1      ====        srai t1, s3, 1
                                                  30'd    4650    : data = 32'h    657C3193    ;    //    sltiu x3 x24 1623      ====        sltiu gp, s8, 1623
                                                  30'd    4651    : data = 32'h    01696BB3    ;    //    or x23 x18 x22      ====        or s7, s2, s6
                                                  30'd    4652    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4653    : data = 32'h    E4D47093    ;    //    andi x1 x8 -435      ====        andi ra, s0, -435
                                                  30'd    4654    : data = 32'h    0C2B7993    ;    //    andi x19 x22 194      ====        andi s3, s6, 194
                                                  30'd    4655    : data = 32'h    00075A93    ;    //    srli x21 x14 0      ====        srli s5, a4, 0
                                                  30'd    4656    : data = 32'h    B7108D13    ;    //    addi x26 x1 -1167      ====        addi s10, ra, -1167
                                                  30'd    4657    : data = 32'h    006A2433    ;    //    slt x8 x20 x6      ====        slt s0, s4, t1
                                                  30'd    4658    : data = 32'h    41595893    ;    //    srai x17 x18 21      ====        srai a7, s2, 21
                                                  30'd    4659    : data = 32'h    B5B5B3B7    ;    //    lui x7 744283      ====        lui t2, 744283
                                                  30'd    4660    : data = 32'h    21B6A993    ;    //    slti x19 x13 539      ====        slti s3, a3, 539
                                                  30'd    4661    : data = 32'h    0E1DA313    ;    //    slti x6 x27 225      ====        slti t1, s11, 225
                                                  30'd    4662    : data = 32'h    87275297    ;    //    auipc x5 553589      ====        auipc t0, 553589
                                                  30'd    4663    : data = 32'h    A7377897    ;    //    auipc x17 684919      ====        auipc a7, 684919
                                                  30'd    4664    : data = 32'h    002D6033    ;    //    or x0 x26 x2      ====        or zero, s10, sp
                                                  30'd    4665    : data = 32'h    01606333    ;    //    or x6 x0 x22      ====        or t1, zero, s6
                                                  30'd    4666    : data = 32'h    7799EF93    ;    //    ori x31 x19 1913      ====        ori t6, s3, 1913
                                                  30'd    4667    : data = 32'h    007CBDB3    ;    //    sltu x27 x25 x7      ====        sltu s11, s9, t2
                                                  30'd    4668    : data = 32'h    51937793    ;    //    andi x15 x6 1305      ====        andi a5, t1, 1305
                                                  30'd    4669    : data = 32'h    410E5333    ;    //    sra x6 x28 x16      ====        sra t1, t3, a6
                                                  30'd    4670    : data = 32'h    40475CB3    ;    //    sra x25 x14 x4      ====        sra s9, a4, tp
                                                  30'd    4671    : data = 32'h    01D6D633    ;    //    srl x12 x13 x29      ====        srl a2, a3, t4
                                                  30'd    4672    : data = 32'h    1AFAA193    ;    //    slti x3 x21 431      ====        slti gp, s5, 431
                                                  30'd    4673    : data = 32'h    9EE62013    ;    //    slti x0 x12 -1554      ====        slti zero, a2, -1554
                                                  30'd    4674    : data = 32'h    B69C4B93    ;    //    xori x23 x24 -1175      ====        xori s7, s8, -1175
                                                  30'd    4675    : data = 32'h    01D2DE13    ;    //    srli x28 x5 29      ====        srli t3, t0, 29
                                                  30'd    4676    : data = 32'h    41365D93    ;    //    srai x27 x12 19      ====        srai s11, a2, 19
                                                  30'd    4677    : data = 32'h    018DC4B3    ;    //    xor x9 x27 x24      ====        xor s1, s11, s8
                                                  30'd    4678    : data = 32'h    00743033    ;    //    sltu x0 x8 x7      ====        sltu zero, s0, t2
                                                  30'd    4679    : data = 32'h    D14BF693    ;    //    andi x13 x23 -748      ====        andi a3, s7, -748
                                                  30'd    4680    : data = 32'h    24FAFC93    ;    //    andi x25 x21 591      ====        andi s9, s5, 591
                                                  30'd    4681    : data = 32'h    00F091B3    ;    //    sll x3 x1 x15      ====        sll gp, ra, a5
                                                  30'd    4682    : data = 32'h    0054B0B3    ;    //    sltu x1 x9 x5      ====        sltu ra, s1, t0
                                                  30'd    4683    : data = 32'h    642CC893    ;    //    xori x17 x25 1602      ====        xori a7, s9, 1602
                                                  30'd    4684    : data = 32'h    013635B3    ;    //    sltu x11 x12 x19      ====        sltu a1, a2, s3
                                                  30'd    4685    : data = 32'h    0124D393    ;    //    srli x7 x9 18      ====        srli t2, s1, 18
                                                  30'd    4686    : data = 32'h    0148D693    ;    //    srli x13 x17 20      ====        srli a3, a7, 20
                                                  30'd    4687    : data = 32'h    40A68EB3    ;    //    sub x29 x13 x10      ====        sub t4, a3, a0
                                                  30'd    4688    : data = 32'h    6107E593    ;    //    ori x11 x15 1552      ====        ori a1, a5, 1552
                                                  30'd    4689    : data = 32'h    8656B013    ;    //    sltiu x0 x13 -1947      ====        sltiu zero, a3, -1947
                                                  30'd    4690    : data = 32'h    01EE22B3    ;    //    slt x5 x28 x30      ====        slt t0, t3, t5
                                                  30'd    4691    : data = 32'h    006B9893    ;    //    slli x17 x23 6      ====        slli a7, s7, 6
                                                  30'd    4692    : data = 32'h    4003D313    ;    //    srai x6 x7 0      ====        srai t1, t2, 0
                                                  30'd    4693    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4694    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4695    : data = 32'h    4111DA13    ;    //    srai x20 x3 17      ====        srai s4, gp, 17
                                                  30'd    4696    : data = 32'h    41358933    ;    //    sub x18 x11 x19      ====        sub s2, a1, s3
                                                  30'd    4697    : data = 32'h    00B6F033    ;    //    and x0 x13 x11      ====        and zero, a3, a1
                                                  30'd    4698    : data = 32'h    00CF17B3    ;    //    sll x15 x30 x12      ====        sll a5, t5, a2
                                                  30'd    4699    : data = 32'h    991A6E17    ;    //    auipc x28 627110      ====        auipc t3, 627110
                                                  30'd    4700    : data = 32'h    00805313    ;    //    srli x6 x0 8      ====        srli t1, zero, 8
                                                  30'd    4701    : data = 32'h    11332A13    ;    //    slti x20 x6 275      ====        slti s4, t1, 275
                                                  30'd    4702    : data = 32'h    0120FAB3    ;    //    and x21 x1 x18      ====        and s5, ra, s2
                                                  30'd    4703    : data = 32'h    007FE833    ;    //    or x16 x31 x7      ====        or a6, t6, t2
                                                  30'd    4704    : data = 32'h    001722B3    ;    //    slt x5 x14 x1      ====        slt t0, a4, ra
                                                  30'd    4705    : data = 32'h    001A86B3    ;    //    add x13 x21 x1      ====        add a3, s5, ra
                                                  30'd    4706    : data = 32'h    63D47B17    ;    //    auipc x22 408903      ====        auipc s6, 408903
                                                  30'd    4707    : data = 32'h    A02BE713    ;    //    ori x14 x23 -1534      ====        ori a4, s7, -1534
                                                  30'd    4708    : data = 32'h    00239A33    ;    //    sll x20 x7 x2      ====        sll s4, t2, sp
                                                  30'd    4709    : data = 32'h    005476B3    ;    //    and x13 x8 x5      ====        and a3, s0, t0
                                                  30'd    4710    : data = 32'h    2FE41417    ;    //    auipc x8 196161      ====        auipc s0, 196161
                                                  30'd    4711    : data = 32'h    4196DFB3    ;    //    sra x31 x13 x25      ====        sra t6, a3, s9
                                                  30'd    4712    : data = 32'h    3C063193    ;    //    sltiu x3 x12 960      ====        sltiu gp, a2, 960
                                                  30'd    4713    : data = 32'h    01644433    ;    //    xor x8 x8 x22      ====        xor s0, s0, s6
                                                  30'd    4714    : data = 32'h    0026DD93    ;    //    srli x27 x13 2      ====        srli s11, a3, 2
                                                  30'd    4715    : data = 32'h    64596993    ;    //    ori x19 x18 1605      ====        ori s3, s2, 1605
                                                  30'd    4716    : data = 32'h    E85BE013    ;    //    ori x0 x23 -379      ====        ori zero, s7, -379
                                                  30'd    4717    : data = 32'h    EBB30713    ;    //    addi x14 x6 -325      ====        addi a4, t1, -325
                                                  30'd    4718    : data = 32'h    A112BE93    ;    //    sltiu x29 x5 -1519      ====        sltiu t4, t0, -1519
                                                  30'd    4719    : data = 32'h    00345813    ;    //    srli x16 x8 3      ====        srli a6, s0, 3
                                                  30'd    4720    : data = 32'h    0BAA8F93    ;    //    addi x31 x21 186      ====        addi t6, s5, 186
                                                  30'd    4721    : data = 32'h    00BB08B3    ;    //    add x17 x22 x11      ====        add a7, s6, a1
                                                  30'd    4722    : data = 32'h    FD65C193    ;    //    xori x3 x11 -42      ====        xori gp, a1, -42
                                                  30'd    4723    : data = 32'h    40F406B3    ;    //    sub x13 x8 x15      ====        sub a3, s0, a5
                                                  30'd    4724    : data = 32'h    F483FB93    ;    //    andi x23 x7 -184      ====        andi s7, t2, -184
                                                  30'd    4725    : data = 32'h    18647193    ;    //    andi x3 x8 390      ====        andi gp, s0, 390
                                                  30'd    4726    : data = 32'h    37172013    ;    //    slti x0 x14 881      ====        slti zero, a4, 881
                                                  30'd    4727    : data = 32'h    003E1E13    ;    //    slli x28 x28 3      ====        slli t3, t3, 3
                                                  30'd    4728    : data = 32'h    40C25633    ;    //    sra x12 x4 x12      ====        sra a2, tp, a2
                                                  30'd    4729    : data = 32'h    404BD433    ;    //    sra x8 x23 x4      ====        sra s0, s7, tp
                                                  30'd    4730    : data = 32'h    014F5293    ;    //    srli x5 x30 20      ====        srli t0, t5, 20
                                                  30'd    4731    : data = 32'h    404153B3    ;    //    sra x7 x2 x4      ====        sra t2, sp, tp
                                                  30'd    4732    : data = 32'h    5E5319B7    ;    //    lui x19 386353      ====        lui s3, 386353
                                                  30'd    4733    : data = 32'h    7F8A0E13    ;    //    addi x28 x20 2040      ====        addi t3, s4, 2040
                                                  30'd    4734    : data = 32'h    400F0733    ;    //    sub x14 x30 x0      ====        sub a4, t5, zero
                                                  30'd    4735    : data = 32'h    01695FB3    ;    //    srl x31 x18 x22      ====        srl t6, s2, s6
                                                  30'd    4736    : data = 32'h    3D7A0E13    ;    //    addi x28 x20 983      ====        addi t3, s4, 983
                                                  30'd    4737    : data = 32'h    0051A9B3    ;    //    slt x19 x3 x5      ====        slt s3, gp, t0
                                                  30'd    4738    : data = 32'h    003929B3    ;    //    slt x19 x18 x3      ====        slt s3, s2, gp
                                                  30'd    4739    : data = 32'h    00790733    ;    //    add x14 x18 x7      ====        add a4, s2, t2
                                                  30'd    4740    : data = 32'h    4FD64113    ;    //    xori x2 x12 1277      ====        xori sp, a2, 1277
                                                  30'd    4741    : data = 32'h    411D8833    ;    //    sub x16 x27 x17      ====        sub a6, s11, a7
                                                  30'd    4742    : data = 32'h    C8662993    ;    //    slti x19 x12 -890      ====        slti s3, a2, -890
                                                  30'd    4743    : data = 32'h    109D7E97    ;    //    auipc x29 68055      ====        auipc t4, 68055
                                                  30'd    4744    : data = 32'h    44DABC93    ;    //    sltiu x25 x21 1101      ====        sltiu s9, s5, 1101
                                                  30'd    4745    : data = 32'h    01841E13    ;    //    slli x28 x8 24      ====        slli t3, s0, 24
                                                  30'd    4746    : data = 32'h    408B5633    ;    //    sra x12 x22 x8      ====        sra a2, s6, s0
                                                  30'd    4747    : data = 32'h    405CDAB3    ;    //    sra x21 x25 x5      ====        sra s5, s9, t0
                                                  30'd    4748    : data = 32'h    00DF2033    ;    //    slt x0 x30 x13      ====        slt zero, t5, a3
                                                  30'd    4749    : data = 32'h    015A8B33    ;    //    add x22 x21 x21      ====        add s6, s5, s5
                                                  30'd    4750    : data = 32'h    01260733    ;    //    add x14 x12 x18      ====        add a4, a2, s2
                                                  30'd    4751    : data = 32'h    03E32113    ;    //    slti x2 x6 62      ====        slti sp, t1, 62
                                                  30'd    4752    : data = 32'h    019FC033    ;    //    xor x0 x31 x25      ====        xor zero, t6, s9
                                                  30'd    4753    : data = 32'h    001A9D33    ;    //    sll x26 x21 x1      ====        sll s10, s5, ra
                                                  30'd    4754    : data = 32'h    41088C33    ;    //    sub x24 x17 x16      ====        sub s8, a7, a6
                                                  30'd    4755    : data = 32'h    0031DE93    ;    //    srli x29 x3 3      ====        srli t4, gp, 3
                                                  30'd    4756    : data = 32'h    004C2FB3    ;    //    slt x31 x24 x4      ====        slt t6, s8, tp
                                                  30'd    4757    : data = 32'h    25C32493    ;    //    slti x9 x6 604      ====        slti s1, t1, 604
                                                  30'd    4758    : data = 32'h    148C0293    ;    //    addi x5 x24 328      ====        addi t0, s8, 328
                                                  30'd    4759    : data = 32'h    00735413    ;    //    srli x8 x6 7      ====        srli s0, t1, 7
                                                  30'd    4760    : data = 32'h    007237B3    ;    //    sltu x15 x4 x7      ====        sltu a5, tp, t2
                                                  30'd    4761    : data = 32'h    56A64493    ;    //    xori x9 x12 1386      ====        xori s1, a2, 1386
                                                  30'd    4762    : data = 32'h    7841FF97    ;    //    auipc x31 492575      ====        auipc t6, 492575
                                                  30'd    4763    : data = 32'h    0036FA33    ;    //    and x20 x13 x3      ====        and s4, a3, gp
                                                  30'd    4764    : data = 32'h    91E2CF93    ;    //    xori x31 x5 -1762      ====        xori t6, t0, -1762
                                                  30'd    4765    : data = 32'h    B1B24793    ;    //    xori x15 x4 -1253      ====        xori a5, tp, -1253
                                                  30'd    4766    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4767    : data = 32'h    010B2733    ;    //    slt x14 x22 x16      ====        slt a4, s6, a6
                                                  30'd    4768    : data = 32'h    01BB1AB3    ;    //    sll x21 x22 x27      ====        sll s5, s6, s11
                                                  30'd    4769    : data = 32'h    00845433    ;    //    srl x8 x8 x8      ====        srl s0, s0, s0
                                                  30'd    4770    : data = 32'h    013EAA33    ;    //    slt x20 x29 x19      ====        slt s4, t4, s3
                                                  30'd    4771    : data = 32'h    5A373193    ;    //    sltiu x3 x14 1443      ====        sltiu gp, a4, 1443
                                                  30'd    4772    : data = 32'h    A7F06E93    ;    //    ori x29 x0 -1409      ====        ori t4, zero, -1409
                                                  30'd    4773    : data = 32'h    01D2D5B3    ;    //    srl x11 x5 x29      ====        srl a1, t0, t4
                                                  30'd    4774    : data = 32'h    014132B3    ;    //    sltu x5 x2 x20      ====        sltu t0, sp, s4
                                                  30'd    4775    : data = 32'h    40708CB3    ;    //    sub x25 x1 x7      ====        sub s9, ra, t2
                                                  30'd    4776    : data = 32'h    01BBECB3    ;    //    or x25 x23 x27      ====        or s9, s7, s11
                                                  30'd    4777    : data = 32'h    010E1DB3    ;    //    sll x27 x28 x16      ====        sll s11, t3, a6
                                                  30'd    4778    : data = 32'h    010FA3B3    ;    //    slt x7 x31 x16      ====        slt t2, t6, a6
                                                  30'd    4779    : data = 32'h    0051ED33    ;    //    or x26 x3 x5      ====        or s10, gp, t0
                                                  30'd    4780    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4781    : data = 32'h    01125AB3    ;    //    srl x21 x4 x17      ====        srl s5, tp, a7
                                                  30'd    4782    : data = 32'h    41EC0FB3    ;    //    sub x31 x24 x30      ====        sub t6, s8, t5
                                                  30'd    4783    : data = 32'h    00A95493    ;    //    srli x9 x18 10      ====        srli s1, s2, 10
                                                  30'd    4784    : data = 32'h    00922EB3    ;    //    slt x29 x4 x9      ====        slt t4, tp, s1
                                                  30'd    4785    : data = 32'h    A599AB13    ;    //    slti x22 x19 -1447      ====        slti s6, s3, -1447
                                                  30'd    4786    : data = 32'h    01A920B3    ;    //    slt x1 x18 x26      ====        slt ra, s2, s10
                                                  30'd    4787    : data = 32'h    F0AC7E93    ;    //    andi x29 x24 -246      ====        andi t4, s8, -246
                                                  30'd    4788    : data = 32'h    00386BB3    ;    //    or x23 x16 x3      ====        or s7, a6, gp
                                                  30'd    4789    : data = 32'h    004F3933    ;    //    sltu x18 x30 x4      ====        sltu s2, t5, tp
                                                  30'd    4790    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4791    : data = 32'h    00814A33    ;    //    xor x20 x2 x8      ====        xor s4, sp, s0
                                                  30'd    4792    : data = 32'h    80940C93    ;    //    addi x25 x8 -2039      ====        addi s9, s0, -2039
                                                  30'd    4793    : data = 32'h    DB6A2C93    ;    //    slti x25 x20 -586      ====        slti s9, s4, -586
                                                  30'd    4794    : data = 32'h    4E19E417    ;    //    auipc x8 319902      ====        auipc s0, 319902
                                                  30'd    4795    : data = 32'h    1C203A93    ;    //    sltiu x21 x0 450      ====        sltiu s5, zero, 450
                                                  30'd    4796    : data = 32'h    4089DE33    ;    //    sra x28 x19 x8      ====        sra t3, s3, s0
                                                  30'd    4797    : data = 32'h    01AD9493    ;    //    slli x9 x27 26      ====        slli s1, s11, 26
                                                  30'd    4798    : data = 32'h    00423133    ;    //    sltu x2 x4 x4      ====        sltu sp, tp, tp
                                                  30'd    4799    : data = 32'h    ADB54013    ;    //    xori x0 x10 -1317      ====        xori zero, a0, -1317
                                                  30'd    4800    : data = 32'h    015681B3    ;    //    add x3 x13 x21      ====        add gp, a3, s5
                                                  30'd    4801    : data = 32'h    BDBEED97    ;    //    auipc x27 777198      ====        auipc s11, 777198
                                                  30'd    4802    : data = 32'h    003BA633    ;    //    slt x12 x23 x3      ====        slt a2, s7, gp
                                                  30'd    4803    : data = 32'h    0149C5B3    ;    //    xor x11 x19 x20      ====        xor a1, s3, s4
                                                  30'd    4804    : data = 32'h    409E52B3    ;    //    sra x5 x28 x9      ====        sra t0, t3, s1
                                                  30'd    4805    : data = 32'h    005A9D13    ;    //    slli x26 x21 5      ====        slli s10, s5, 5
                                                  30'd    4806    : data = 32'h    017C0733    ;    //    add x14 x24 x23      ====        add a4, s8, s7
                                                  30'd    4807    : data = 32'h    00C27633    ;    //    and x12 x4 x12      ====        and a2, tp, a2
                                                  30'd    4808    : data = 32'h    3B426017    ;    //    auipc x0 242726      ====        auipc zero, 242726
                                                  30'd    4809    : data = 32'h    81D2BF93    ;    //    sltiu x31 x5 -2019      ====        sltiu t6, t0, -2019
                                                  30'd    4810    : data = 32'h    014B23B3    ;    //    slt x7 x22 x20      ====        slt t2, s6, s4
                                                  30'd    4811    : data = 32'h    411AD2B3    ;    //    sra x5 x21 x17      ====        sra t0, s5, a7
                                                  30'd    4812    : data = 32'h    AE30BD13    ;    //    sltiu x26 x1 -1309      ====        sltiu s10, ra, -1309
                                                  30'd    4813    : data = 32'h    8259E393    ;    //    ori x7 x19 -2011      ====        ori t2, s3, -2011
                                                  30'd    4814    : data = 32'h    2472F493    ;    //    andi x9 x5 583      ====        andi s1, t0, 583
                                                  30'd    4815    : data = 32'h    01CB9613    ;    //    slli x12 x23 28      ====        slli a2, s7, 28
                                                  30'd    4816    : data = 32'h    9F2EEB93    ;    //    ori x23 x29 -1550      ====        ori s7, t4, -1550
                                                  30'd    4817    : data = 32'h    18310A13    ;    //    addi x20 x2 387      ====        addi s4, sp, 387
                                                  30'd    4818    : data = 32'h    4054D6B3    ;    //    sra x13 x9 x5      ====        sra a3, s1, t0
                                                  30'd    4819    : data = 32'h    749AF797    ;    //    auipc x15 477615      ====        auipc a5, 477615
                                                  30'd    4820    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4821    : data = 32'h    5D076713    ;    //    ori x14 x14 1488      ====        ori a4, a4, 1488
                                                  30'd    4822    : data = 32'h    0018E6B3    ;    //    or x13 x17 x1      ====        or a3, a7, ra
                                                  30'd    4823    : data = 32'h    019E1DB3    ;    //    sll x27 x28 x25      ====        sll s11, t3, s9
                                                  30'd    4824    : data = 32'h    000B33B3    ;    //    sltu x7 x22 x0      ====        sltu t2, s6, zero
                                                  30'd    4825    : data = 32'h    016E29B3    ;    //    slt x19 x28 x22      ====        slt s3, t3, s6
                                                  30'd    4826    : data = 32'h    9D0B3813    ;    //    sltiu x16 x22 -1584      ====        sltiu a6, s6, -1584
                                                  30'd    4827    : data = 32'h    31A78293    ;    //    addi x5 x15 794      ====        addi t0, a5, 794
                                                  30'd    4828    : data = 32'h    01E14333    ;    //    xor x6 x2 x30      ====        xor t1, sp, t5
                                                  30'd    4829    : data = 32'h    40E18733    ;    //    sub x14 x3 x14      ====        sub a4, gp, a4
                                                  30'd    4830    : data = 32'h    63F5B997    ;    //    auipc x19 409435      ====        auipc s3, 409435
                                                  30'd    4831    : data = 32'h    D7314713    ;    //    xori x14 x2 -653      ====        xori a4, sp, -653
                                                  30'd    4832    : data = 32'h    01936033    ;    //    or x0 x6 x25      ====        or zero, t1, s9
                                                  30'd    4833    : data = 32'h    00D8EB33    ;    //    or x22 x17 x13      ====        or s6, a7, a3
                                                  30'd    4834    : data = 32'h    75B76717    ;    //    auipc x14 482166      ====        auipc a4, 482166
                                                  30'd    4835    : data = 32'h    00609093    ;    //    slli x1 x1 6      ====        slli ra, ra, 6
                                                  30'd    4836    : data = 32'h    D4233F93    ;    //    sltiu x31 x6 -702      ====        sltiu t6, t1, -702
                                                  30'd    4837    : data = 32'h    471D1317    ;    //    auipc x6 291281      ====        auipc t1, 291281
                                                  30'd    4838    : data = 32'h    4086D693    ;    //    srai x13 x13 8      ====        srai a3, a3, 8
                                                  30'd    4839    : data = 32'h    003C2133    ;    //    slt x2 x24 x3      ====        slt sp, s8, gp
                                                  30'd    4840    : data = 32'h    41495C33    ;    //    sra x24 x18 x20      ====        sra s8, s2, s4
                                                  30'd    4841    : data = 32'h    C486F793    ;    //    andi x15 x13 -952      ====        andi a5, a3, -952
                                                  30'd    4842    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4843    : data = 32'h    005F64B3    ;    //    or x9 x30 x5      ====        or s1, t5, t0
                                                  30'd    4844    : data = 32'h    00DF47B3    ;    //    xor x15 x30 x13      ====        xor a5, t5, a3
                                                  30'd    4845    : data = 32'h    5E31EB93    ;    //    ori x23 x3 1507      ====        ori s7, gp, 1507
                                                  30'd    4846    : data = 32'h    01EF5293    ;    //    srli x5 x30 30      ====        srli t0, t5, 30
                                                  30'd    4847    : data = 32'h    01D11D33    ;    //    sll x26 x2 x29      ====        sll s10, sp, t4
                                                  30'd    4848    : data = 32'h    01D6E5B3    ;    //    or x11 x13 x29      ====        or a1, a3, t4
                                                  30'd    4849    : data = 32'h    401CDB93    ;    //    srai x23 x25 1      ====        srai s7, s9, 1
                                                  30'd    4850    : data = 32'h    63E56613    ;    //    ori x12 x10 1598      ====        ori a2, a0, 1598
                                                  30'd    4851    : data = 32'h    011747B3    ;    //    xor x15 x14 x17      ====        xor a5, a4, a7
                                                  30'd    4852    : data = 32'h    000E58B3    ;    //    srl x17 x28 x0      ====        srl a7, t3, zero
                                                  30'd    4853    : data = 32'h    000B4D33    ;    //    xor x26 x22 x0      ====        xor s10, s6, zero
                                                  30'd    4854    : data = 32'h    84EB2913    ;    //    slti x18 x22 -1970      ====        slti s2, s6, -1970
                                                  30'd    4855    : data = 32'h    015F5DB3    ;    //    srl x27 x30 x21      ====        srl s11, t5, s5
                                                  30'd    4856    : data = 32'h    007ADC93    ;    //    srli x25 x21 7      ====        srli s9, s5, 7
                                                  30'd    4857    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4858    : data = 32'h    417C5E33    ;    //    sra x28 x24 x23      ====        sra t3, s8, s7
                                                  30'd    4859    : data = 32'h    002123B3    ;    //    slt x7 x2 x2      ====        slt t2, sp, sp
                                                  30'd    4860    : data = 32'h    9C96A897    ;    //    auipc x17 641386      ====        auipc a7, 641386
                                                  30'd    4861    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4862    : data = 32'h    011E9B93    ;    //    slli x23 x29 17      ====        slli s7, t4, 17
                                                  30'd    4863    : data = 32'h    01CFF9B3    ;    //    and x19 x31 x28      ====        and s3, t6, t3
                                                  30'd    4864    : data = 32'h    000CADB3    ;    //    slt x27 x25 x0      ====        slt s11, s9, zero
                                                  30'd    4865    : data = 32'h    0120BB33    ;    //    sltu x22 x1 x18      ====        sltu s6, ra, s2
                                                  30'd    4866    : data = 32'h    E444FE13    ;    //    andi x28 x9 -444      ====        andi t3, s1, -444
                                                  30'd    4867    : data = 32'h    01CCDEB3    ;    //    srl x29 x25 x28      ====        srl t4, s9, t3
                                                  30'd    4868    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4869    : data = 32'h    404C5A93    ;    //    srai x21 x24 4      ====        srai s5, s8, 4
                                                  30'd    4870    : data = 32'h    01739E93    ;    //    slli x29 x7 23      ====        slli t4, t2, 23
                                                  30'd    4871    : data = 32'h    40BF54B3    ;    //    sra x9 x30 x11      ====        sra s1, t5, a1
                                                  30'd    4872    : data = 32'h    0189BA33    ;    //    sltu x20 x19 x24      ====        sltu s4, s3, s8
                                                  30'd    4873    : data = 32'h    0025C733    ;    //    xor x14 x11 x2      ====        xor a4, a1, sp
                                                  30'd    4874    : data = 32'h    41AB03B3    ;    //    sub x7 x22 x26      ====        sub t2, s6, s10
                                                  30'd    4875    : data = 32'h    00D35913    ;    //    srli x18 x6 13      ====        srli s2, t1, 13
                                                  30'd    4876    : data = 32'h    0179EEB3    ;    //    or x29 x19 x23      ====        or t4, s3, s7
                                                  30'd    4877    : data = 32'h    012730B3    ;    //    sltu x1 x14 x18      ====        sltu ra, a4, s2
                                                  30'd    4878    : data = 32'h    0077CB33    ;    //    xor x22 x15 x7      ====        xor s6, a5, t2
                                                  30'd    4879    : data = 32'h    006A3E33    ;    //    sltu x28 x20 x6      ====        sltu t3, s4, t1
                                                  30'd    4880    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4881    : data = 32'h    009A08B3    ;    //    add x17 x20 x9      ====        add a7, s4, s1
                                                  30'd    4882    : data = 32'h    01419133    ;    //    sll x2 x3 x20      ====        sll sp, gp, s4
                                                  30'd    4883    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4884    : data = 32'h    AAE00593    ;    //    addi x11 x0 -1362      ====        addi a1, zero, -1362
                                                  30'd    4885    : data = 32'h    FFBA7693    ;    //    andi x13 x20 -5      ====        andi a3, s4, -5
                                                  30'd    4886    : data = 32'h    06436B93    ;    //    ori x23 x6 100      ====        ori s7, t1, 100
                                                  30'd    4887    : data = 32'h    41EEDC13    ;    //    srai x24 x29 30      ====        srai s8, t4, 30
                                                  30'd    4888    : data = 32'h    007469B3    ;    //    or x19 x8 x7      ====        or s3, s0, t2
                                                  30'd    4889    : data = 32'h    3BD7B613    ;    //    sltiu x12 x15 957      ====        sltiu a2, a5, 957
                                                  30'd    4890    : data = 32'h    00B2BD33    ;    //    sltu x26 x5 x11      ====        sltu s10, t0, a1
                                                  30'd    4891    : data = 32'h    0183D013    ;    //    srli x0 x7 24      ====        srli zero, t2, 24
                                                  30'd    4892    : data = 32'h    8BD16013    ;    //    ori x0 x2 -1859      ====        ori zero, sp, -1859
                                                  30'd    4893    : data = 32'h    97DEA713    ;    //    slti x14 x29 -1667      ====        slti a4, t4, -1667
                                                  30'd    4894    : data = 32'h    00DD3D33    ;    //    sltu x26 x26 x13      ====        sltu s10, s10, a3
                                                  30'd    4895    : data = 32'h    01D79F93    ;    //    slli x31 x15 29      ====        slli t6, a5, 29
                                                  30'd    4896    : data = 32'h    41E25C93    ;    //    srai x25 x4 30      ====        srai s9, tp, 30
                                                  30'd    4897    : data = 32'h    01AF2633    ;    //    slt x12 x30 x26      ====        slt a2, t5, s10
                                                  30'd    4898    : data = 32'h    40295D93    ;    //    srai x27 x18 2      ====        srai s11, s2, 2
                                                  30'd    4899    : data = 32'h    4085D693    ;    //    srai x13 x11 8      ====        srai a3, a1, 8
                                                  30'd    4900    : data = 32'h    01174DB3    ;    //    xor x27 x14 x17      ====        xor s11, a4, a7
                                                  30'd    4901    : data = 32'h    A032A793    ;    //    slti x15 x5 -1533      ====        slti a5, t0, -1533
                                                  30'd    4902    : data = 32'h    AC80C017    ;    //    auipc x0 706572      ====        auipc zero, 706572
                                                  30'd    4903    : data = 32'h    12F77D93    ;    //    andi x27 x14 303      ====        andi s11, a4, 303
                                                  30'd    4904    : data = 32'h    001B78B3    ;    //    and x17 x22 x1      ====        and a7, s6, ra
                                                  30'd    4905    : data = 32'h    001DBCB3    ;    //    sltu x25 x27 x1      ====        sltu s9, s11, ra
                                                  30'd    4906    : data = 32'h    0036FDB3    ;    //    and x27 x13 x3      ====        and s11, a3, gp
                                                  30'd    4907    : data = 32'h    006DAFB3    ;    //    slt x31 x27 x6      ====        slt t6, s11, t1
                                                  30'd    4908    : data = 32'h    57437413    ;    //    andi x8 x6 1396      ====        andi s0, t1, 1396
                                                  30'd    4909    : data = 32'h    012949B3    ;    //    xor x19 x18 x18      ====        xor s3, s2, s2
                                                  30'd    4910    : data = 32'h    0001D293    ;    //    srli x5 x3 0      ====        srli t0, gp, 0
                                                  30'd    4911    : data = 32'h    00D69B33    ;    //    sll x22 x13 x13      ====        sll s6, a3, a3
                                                  30'd    4912    : data = 32'h    79788B93    ;    //    addi x23 x17 1943      ====        addi s7, a7, 1943
                                                  30'd    4913    : data = 32'h    41995493    ;    //    srai x9 x18 25      ====        srai s1, s2, 25
                                                  30'd    4914    : data = 32'h    6E4FAE13    ;    //    slti x28 x31 1764      ====        slti t3, t6, 1764
                                                  30'd    4915    : data = 32'h    4149DB93    ;    //    srai x23 x19 20      ====        srai s7, s3, 20
                                                  30'd    4916    : data = 32'h    01405D93    ;    //    srli x27 x0 20      ====        srli s11, zero, 20
                                                  30'd    4917    : data = 32'h    01728D33    ;    //    add x26 x5 x23      ====        add s10, t0, s7
                                                  30'd    4918    : data = 32'h    01C45E93    ;    //    srli x29 x8 28      ====        srli t4, s0, 28
                                                  30'd    4919    : data = 32'h    00B6BE33    ;    //    sltu x28 x13 x11      ====        sltu t3, a3, a1
                                                  30'd    4920    : data = 32'h    B46AB993    ;    //    sltiu x19 x21 -1210      ====        sltiu s3, s5, -1210
                                                  30'd    4921    : data = 32'h    0002DA93    ;    //    srli x21 x5 0      ====        srli s5, t0, 0
                                                  30'd    4922    : data = 32'h    40D15433    ;    //    sra x8 x2 x13      ====        sra s0, sp, a3
                                                  30'd    4923    : data = 32'h    015993B3    ;    //    sll x7 x19 x21      ====        sll t2, s3, s5
                                                  30'd    4924    : data = 32'h    01BDDD13    ;    //    srli x26 x27 27      ====        srli s10, s11, 27
                                                  30'd    4925    : data = 32'h    00ED3333    ;    //    sltu x6 x26 x14      ====        sltu t1, s10, a4
                                                  30'd    4926    : data = 32'h    007F7633    ;    //    and x12 x30 x7      ====        and a2, t5, t2
                                                  30'd    4927    : data = 32'h    0036D2B3    ;    //    srl x5 x13 x3      ====        srl t0, a3, gp
                                                  30'd    4928    : data = 32'h    D08CF393    ;    //    andi x7 x25 -760      ====        andi t2, s9, -760
                                                  30'd    4929    : data = 32'h    20E8E293    ;    //    ori x5 x17 526      ====        ori t0, a7, 526
                                                  30'd    4930    : data = 32'h    01361A93    ;    //    slli x21 x12 19      ====        slli s5, a2, 19
                                                  30'd    4931    : data = 32'h    B138A093    ;    //    slti x1 x17 -1261      ====        slti ra, a7, -1261
                                                  30'd    4932    : data = 32'h    405A06B3    ;    //    sub x13 x20 x5      ====        sub a3, s4, t0
                                                  30'd    4933    : data = 32'h    ED658B13    ;    //    addi x22 x11 -298      ====        addi s6, a1, -298
                                                  30'd    4934    : data = 32'h    41FE86B3    ;    //    sub x13 x29 x31      ====        sub a3, t4, t6
                                                  30'd    4935    : data = 32'h    01C441B3    ;    //    xor x3 x8 x28      ====        xor gp, s0, t3
                                                  30'd    4936    : data = 32'h    0012C6B3    ;    //    xor x13 x5 x1      ====        xor a3, t0, ra
                                                  30'd    4937    : data = 32'h    01DC1933    ;    //    sll x18 x24 x29      ====        sll s2, s8, t4
                                                  30'd    4938    : data = 32'h    4176D793    ;    //    srai x15 x13 23      ====        srai a5, a3, 23
                                                  30'd    4939    : data = 32'h    01662BB3    ;    //    slt x23 x12 x22      ====        slt s7, a2, s6
                                                  30'd    4940    : data = 32'h    41775C33    ;    //    sra x24 x14 x23      ====        sra s8, a4, s7
                                                  30'd    4941    : data = 32'h    E3FA4313    ;    //    xori x6 x20 -449      ====        xori t1, s4, -449
                                                  30'd    4942    : data = 32'h    01448433    ;    //    add x8 x9 x20      ====        add s0, s1, s4
                                                  30'd    4943    : data = 32'h    01CF80B3    ;    //    add x1 x31 x28      ====        add ra, t6, t3
                                                  30'd    4944    : data = 32'h    01EAD333    ;    //    srl x6 x21 x30      ====        srl t1, s5, t5
                                                  30'd    4945    : data = 32'h    0087BE33    ;    //    sltu x28 x15 x8      ====        sltu t3, a5, s0
                                                  30'd    4946    : data = 32'h    0030CEB3    ;    //    xor x29 x1 x3      ====        xor t4, ra, gp
                                                  30'd    4947    : data = 32'h    000F9993    ;    //    slli x19 x31 0      ====        slli s3, t6, 0
                                                  30'd    4948    : data = 32'h    F765B593    ;    //    sltiu x11 x11 -138      ====        sltiu a1, a1, -138
                                                  30'd    4949    : data = 32'h    41BA81B3    ;    //    sub x3 x21 x27      ====        sub gp, s5, s11
                                                  30'd    4950    : data = 32'h    417B86B3    ;    //    sub x13 x23 x23      ====        sub a3, s7, s7
                                                  30'd    4951    : data = 32'h    1045E697    ;    //    auipc x13 66654      ====        auipc a3, 66654
                                                  30'd    4952    : data = 32'h    40C257B3    ;    //    sra x15 x4 x12      ====        sra a5, tp, a2
                                                  30'd    4953    : data = 32'h    014A2AB3    ;    //    slt x21 x20 x20      ====        slt s5, s4, s4
                                                  30'd    4954    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4955    : data = 32'h    41B584B3    ;    //    sub x9 x11 x27      ====        sub s1, a1, s11
                                                  30'd    4956    : data = 32'h    4013DC33    ;    //    sra x24 x7 x1      ====        sra s8, t2, ra
                                                  30'd    4957    : data = 32'h    2472E393    ;    //    ori x7 x5 583      ====        ori t2, t0, 583
                                                  30'd    4958    : data = 32'h    5A4DAA93    ;    //    slti x21 x27 1444      ====        slti s5, s11, 1444
                                                  30'd    4959    : data = 32'h    AA2C8713    ;    //    addi x14 x25 -1374      ====        addi a4, s9, -1374
                                                  30'd    4960    : data = 32'h    41B8D6B3    ;    //    sra x13 x17 x27      ====        sra a3, a7, s11
                                                  30'd    4961    : data = 32'h    6A8D3F97    ;    //    auipc x31 436435      ====        auipc t6, 436435
                                                  30'd    4962    : data = 32'h    40D407B3    ;    //    sub x15 x8 x13      ====        sub a5, s0, a3
                                                  30'd    4963    : data = 32'h    01AC1293    ;    //    slli x5 x24 26      ====        slli t0, s8, 26
                                                  30'd    4964    : data = 32'h    91AD4F93    ;    //    xori x31 x26 -1766      ====        xori t6, s10, -1766
                                                  30'd    4965    : data = 32'h    010ED633    ;    //    srl x12 x29 x16      ====        srl a2, t4, a6
                                                  30'd    4966    : data = 32'h    00B7BCB3    ;    //    sltu x25 x15 x11      ====        sltu s9, a5, a1
                                                  30'd    4967    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4968    : data = 32'h    41F84B93    ;    //    xori x23 x16 1055      ====        xori s7, a6, 1055
                                                  30'd    4969    : data = 32'h    A2F6F713    ;    //    andi x14 x13 -1489      ====        andi a4, a3, -1489
                                                  30'd    4970    : data = 32'h    ED3ADE37    ;    //    lui x28 971693      ====        lui t3, 971693
                                                  30'd    4971    : data = 32'h    00FE0C33    ;    //    add x24 x28 x15      ====        add s8, t3, a5
                                                  30'd    4972    : data = 32'h    07560113    ;    //    addi x2 x12 117      ====        addi sp, a2, 117
                                                  30'd    4973    : data = 32'h    400B0333    ;    //    sub x6 x22 x0      ====        sub t1, s6, zero
                                                  30'd    4974    : data = 32'h    50BFF693    ;    //    andi x13 x31 1291      ====        andi a3, t6, 1291
                                                  30'd    4975    : data = 32'h    01CAC5B3    ;    //    xor x11 x21 x28      ====        xor a1, s5, t3
                                                  30'd    4976    : data = 32'h    41425113    ;    //    srai x2 x4 20      ====        srai sp, tp, 20
                                                  30'd    4977    : data = 32'h    1DF491B7    ;    //    lui x3 122697      ====        lui gp, 122697
                                                  30'd    4978    : data = 32'h    0027C593    ;    //    xori x11 x15 2      ====        xori a1, a5, 2
                                                  30'd    4979    : data = 32'h    411855B3    ;    //    sra x11 x16 x17      ====        sra a1, a6, a7
                                                  30'd    4980    : data = 32'h    0050B333    ;    //    sltu x6 x1 x5      ====        sltu t1, ra, t0
                                                  30'd    4981    : data = 32'h    67AC7C93    ;    //    andi x25 x24 1658      ====        andi s9, s8, 1658
                                                  30'd    4982    : data = 32'h    0063DDB3    ;    //    srl x27 x7 x6      ====        srl s11, t2, t1
                                                  30'd    4983    : data = 32'h    019482B3    ;    //    add x5 x9 x25      ====        add t0, s1, s9
                                                  30'd    4984    : data = 32'h    41CDD2B3    ;    //    sra x5 x27 x28      ====        sra t0, s11, t3
                                                  30'd    4985    : data = 32'h    00B23333    ;    //    sltu x6 x4 x11      ====        sltu t1, tp, a1
                                                  30'd    4986    : data = 32'h    0014E8B3    ;    //    or x17 x9 x1      ====        or a7, s1, ra
                                                  30'd    4987    : data = 32'h    407B5A93    ;    //    srai x21 x22 7      ====        srai s5, s6, 7
                                                  30'd    4988    : data = 32'h    01536A33    ;    //    or x20 x6 x21      ====        or s4, t1, s5
                                                  30'd    4989    : data = 32'h    DE066637    ;    //    lui x12 909414      ====        lui a2, 909414
                                                  30'd    4990    : data = 32'h    40455593    ;    //    srai x11 x10 4      ====        srai a1, a0, 4
                                                  30'd    4991    : data = 32'h    00DBE9B3    ;    //    or x19 x23 x13      ====        or s3, s7, a3
                                                  30'd    4992    : data = 32'h    015AB033    ;    //    sltu x0 x21 x21      ====        sltu zero, s5, s5
                                                  30'd    4993    : data = 32'h    315EF993    ;    //    andi x19 x29 789      ====        andi s3, t4, 789
                                                  30'd    4994    : data = 32'h    BCB97E13    ;    //    andi x28 x18 -1077      ====        andi t3, s2, -1077
                                                  30'd    4995    : data = 32'h    41A00AB3    ;    //    sub x21 x0 x26      ====        sub s5, zero, s10
                                                  30'd    4996    : data = 32'h    005C5293    ;    //    srli x5 x24 5      ====        srli t0, s8, 5
                                                  30'd    4997    : data = 32'h    017D1FB3    ;    //    sll x31 x26 x23      ====        sll t6, s10, s7
                                                  30'd    4998    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    4999    : data = 32'h    A37DBE93    ;    //    sltiu x29 x27 -1481      ====        sltiu t4, s11, -1481
                                                  30'd    5000    : data = 32'h    01E6B4B3    ;    //    sltu x9 x13 x30      ====        sltu s1, a3, t5
                                                  30'd    5001    : data = 32'h    11C3FB13    ;    //    andi x22 x7 284      ====        andi s6, t2, 284
                                                  30'd    5002    : data = 32'h    01957633    ;    //    and x12 x10 x25      ====        and a2, a0, s9
                                                  30'd    5003    : data = 32'h    01EEFEB3    ;    //    and x29 x29 x30      ====        and t4, t4, t5
                                                  30'd    5004    : data = 32'h    0143A2B3    ;    //    slt x5 x7 x20      ====        slt t0, t2, s4
                                                  30'd    5005    : data = 32'h    007DDA33    ;    //    srl x20 x27 x7      ====        srl s4, s11, t2
                                                  30'd    5006    : data = 32'h    C8902DB7    ;    //    lui x27 821506      ====        lui s11, 821506
                                                  30'd    5007    : data = 32'h    8B47A493    ;    //    slti x9 x15 -1868      ====        slti s1, a5, -1868
                                                  30'd    5008    : data = 32'h    00D88433    ;    //    add x8 x17 x13      ====        add s0, a7, a3
                                                  30'd    5009    : data = 32'h    00B98433    ;    //    add x8 x19 x11      ====        add s0, s3, a1
                                                  30'd    5010    : data = 32'h    004451B3    ;    //    srl x3 x8 x4      ====        srl gp, s0, tp
                                                  30'd    5011    : data = 32'h    00E95D93    ;    //    srli x27 x18 14      ====        srli s11, s2, 14
                                                  30'd    5012    : data = 32'h    00C09C13    ;    //    slli x24 x1 12      ====        slli s8, ra, 12
                                                  30'd    5013    : data = 32'h    B8F3A617    ;    //    auipc x12 757562      ====        auipc a2, 757562
                                                  30'd    5014    : data = 32'h    00E77933    ;    //    and x18 x14 x14      ====        and s2, a4, a4
                                                  30'd    5015    : data = 32'h    000231B3    ;    //    sltu x3 x4 x0      ====        sltu gp, tp, zero
                                                  30'd    5016    : data = 32'h    00F75433    ;    //    srl x8 x14 x15      ====        srl s0, a4, a5
                                                  30'd    5017    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5018    : data = 32'h    012053B3    ;    //    srl x7 x0 x18      ====        srl t2, zero, s2
                                                  30'd    5019    : data = 32'h    012C9A13    ;    //    slli x20 x25 18      ====        slli s4, s9, 18
                                                  30'd    5020    : data = 32'h    41C859B3    ;    //    sra x19 x16 x28      ====        sra s3, a6, t3
                                                  30'd    5021    : data = 32'h    A32E6013    ;    //    ori x0 x28 -1486      ====        ori zero, t3, -1486
                                                  30'd    5022    : data = 32'h    009ED7B3    ;    //    srl x15 x29 x9      ====        srl a5, t4, s1
                                                  30'd    5023    : data = 32'h    7AA0C993    ;    //    xori x19 x1 1962      ====        xori s3, ra, 1962
                                                  30'd    5024    : data = 32'h    01195E93    ;    //    srli x29 x18 17      ====        srli t4, s2, 17
                                                  30'd    5025    : data = 32'h    11ED5797    ;    //    auipc x15 73429      ====        auipc a5, 73429
                                                  30'd    5026    : data = 32'h    419188B3    ;    //    sub x17 x3 x25      ====        sub a7, gp, s9
                                                  30'd    5027    : data = 32'h    011A0C33    ;    //    add x24 x20 x17      ====        add s8, s4, a7
                                                  30'd    5028    : data = 32'h    006A6C33    ;    //    or x24 x20 x6      ====        or s8, s4, t1
                                                  30'd    5029    : data = 32'h    5200F613    ;    //    andi x12 x1 1312      ====        andi a2, ra, 1312
                                                  30'd    5030    : data = 32'h    00185613    ;    //    srli x12 x16 1      ====        srli a2, a6, 1
                                                  30'd    5031    : data = 32'h    00601833    ;    //    sll x16 x0 x6      ====        sll a6, zero, t1
                                                  30'd    5032    : data = 32'h    00BB0BB3    ;    //    add x23 x22 x11      ====        add s7, s6, a1
                                                  30'd    5033    : data = 32'h    008E5713    ;    //    srli x14 x28 8      ====        srli a4, t3, 8
                                                  30'd    5034    : data = 32'h    1C430B13    ;    //    addi x22 x6 452      ====        addi s6, t1, 452
                                                  30'd    5035    : data = 32'h    00335E13    ;    //    srli x28 x6 3      ====        srli t3, t1, 3
                                                  30'd    5036    : data = 32'h    01EAEBB3    ;    //    or x23 x21 x30      ====        or s7, s5, t5
                                                  30'd    5037    : data = 32'h    6A2DC093    ;    //    xori x1 x27 1698      ====        xori ra, s11, 1698
                                                  30'd    5038    : data = 32'h    11F67613    ;    //    andi x12 x12 287      ====        andi a2, a2, 287
                                                  30'd    5039    : data = 32'h    00B21593    ;    //    slli x11 x4 11      ====        slli a1, tp, 11
                                                  30'd    5040    : data = 32'h    E8673393    ;    //    sltiu x7 x14 -378      ====        sltiu t2, a4, -378
                                                  30'd    5041    : data = 32'h    00653EB3    ;    //    sltu x29 x10 x6      ====        sltu t4, a0, t1
                                                  30'd    5042    : data = 32'h    003E0733    ;    //    add x14 x28 x3      ====        add a4, t3, gp
                                                  30'd    5043    : data = 32'h    001C1B33    ;    //    sll x22 x24 x1      ====        sll s6, s8, ra
                                                  30'd    5044    : data = 32'h    EA2C2297    ;    //    auipc x5 959170      ====        auipc t0, 959170
                                                  30'd    5045    : data = 32'h    01DE86B3    ;    //    add x13 x29 x29      ====        add a3, t4, t4
                                                  30'd    5046    : data = 32'h    01D8ADB3    ;    //    slt x27 x17 x29      ====        slt s11, a7, t4
                                                  30'd    5047    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5048    : data = 32'h    0059D0B3    ;    //    srl x1 x19 x5      ====        srl ra, s3, t0
                                                  30'd    5049    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5050    : data = 32'h    00624433    ;    //    xor x8 x4 x6      ====        xor s0, tp, t1
                                                  30'd    5051    : data = 32'h    00585713    ;    //    srli x14 x16 5      ====        srli a4, a6, 5
                                                  30'd    5052    : data = 32'h    013286B3    ;    //    add x13 x5 x19      ====        add a3, t0, s3
                                                  30'd    5053    : data = 32'h    40515C93    ;    //    srai x25 x2 5      ====        srai s9, sp, 5
                                                  30'd    5054    : data = 32'h    41770AB3    ;    //    sub x21 x14 x23      ====        sub s5, a4, s7
                                                  30'd    5055    : data = 32'h    40A756B3    ;    //    sra x13 x14 x10      ====        sra a3, a4, a0
                                                  30'd    5056    : data = 32'h    40B9DA13    ;    //    srai x20 x19 11      ====        srai s4, s3, 11
                                                  30'd    5057    : data = 32'h    EAA48613    ;    //    addi x12 x9 -342      ====        addi a2, s1, -342
                                                  30'd    5058    : data = 32'h    00F9AE33    ;    //    slt x28 x19 x15      ====        slt t3, s3, a5
                                                  30'd    5059    : data = 32'h    40D90CB3    ;    //    sub x25 x18 x13      ====        sub s9, s2, a3
                                                  30'd    5060    : data = 32'h    DF70A693    ;    //    slti x13 x1 -521      ====        slti a3, ra, -521
                                                  30'd    5061    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5062    : data = 32'h    38BB4B13    ;    //    xori x22 x22 907      ====        xori s6, s6, 907
                                                  30'd    5063    : data = 32'h    E23DA5B7    ;    //    lui x11 926682      ====        lui a1, 926682
                                                  30'd    5064    : data = 32'h    00919633    ;    //    sll x12 x3 x9      ====        sll a2, gp, s1
                                                  30'd    5065    : data = 32'h    41AD8133    ;    //    sub x2 x27 x26      ====        sub sp, s11, s10
                                                  30'd    5066    : data = 32'h    78F61D37    ;    //    lui x26 495457      ====        lui s10, 495457
                                                  30'd    5067    : data = 32'h    42432597    ;    //    auipc x11 271410      ====        auipc a1, 271410
                                                  30'd    5068    : data = 32'h    00672FB3    ;    //    slt x31 x14 x6      ====        slt t6, a4, t1
                                                  30'd    5069    : data = 32'h    51A50097    ;    //    auipc x1 334416      ====        auipc ra, 334416
                                                  30'd    5070    : data = 32'h    EA6D6113    ;    //    ori x2 x26 -346      ====        ori sp, s10, -346
                                                  30'd    5071    : data = 32'h    8EC98193    ;    //    addi x3 x19 -1812      ====        addi gp, s3, -1812
                                                  30'd    5072    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5073    : data = 32'h    C1EAB013    ;    //    sltiu x0 x21 -994      ====        sltiu zero, s5, -994
                                                  30'd    5074    : data = 32'h    0135FB33    ;    //    and x22 x11 x19      ====        and s6, a1, s3
                                                  30'd    5075    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5076    : data = 32'h    003841B3    ;    //    xor x3 x16 x3      ====        xor gp, a6, gp
                                                  30'd    5077    : data = 32'h    41DD5D33    ;    //    sra x26 x26 x29      ====        sra s10, s10, t4
                                                  30'd    5078    : data = 32'h    DEB3E793    ;    //    ori x15 x7 -533      ====        ori a5, t2, -533
                                                  30'd    5079    : data = 32'h    003335B3    ;    //    sltu x11 x6 x3      ====        sltu a1, t1, gp
                                                  30'd    5080    : data = 32'h    40275693    ;    //    srai x13 x14 2      ====        srai a3, a4, 2
                                                  30'd    5081    : data = 32'h    00396D33    ;    //    or x26 x18 x3      ====        or s10, s2, gp
                                                  30'd    5082    : data = 32'h    01F58133    ;    //    add x2 x11 x31      ====        add sp, a1, t6
                                                  30'd    5083    : data = 32'h    9DE8AA13    ;    //    slti x20 x17 -1570      ====        slti s4, a7, -1570
                                                  30'd    5084    : data = 32'h    017F1F93    ;    //    slli x31 x30 23      ====        slli t6, t5, 23
                                                  30'd    5085    : data = 32'h    C4A860B7    ;    //    lui x1 805510      ====        lui ra, 805510
                                                  30'd    5086    : data = 32'h    017C3EB3    ;    //    sltu x29 x24 x23      ====        sltu t4, s8, s7
                                                  30'd    5087    : data = 32'h    000953B3    ;    //    srl x7 x18 x0      ====        srl t2, s2, zero
                                                  30'd    5088    : data = 32'h    00935393    ;    //    srli x7 x6 9      ====        srli t2, t1, 9
                                                  30'd    5089    : data = 32'h    01759B93    ;    //    slli x23 x11 23      ====        slli s7, a1, 23
                                                  30'd    5090    : data = 32'h    27EB2393    ;    //    slti x7 x22 638      ====        slti t2, s6, 638
                                                  30'd    5091    : data = 32'h    A451F913    ;    //    andi x18 x3 -1467      ====        andi s2, gp, -1467
                                                  30'd    5092    : data = 32'h    40F7D8B3    ;    //    sra x17 x15 x15      ====        sra a7, a5, a5
                                                  30'd    5093    : data = 32'h    4132DE13    ;    //    srai x28 x5 19      ====        srai t3, t0, 19
                                                  30'd    5094    : data = 32'h    93898413    ;    //    addi x8 x19 -1736      ====        addi s0, s3, -1736
                                                  30'd    5095    : data = 32'h    D3BBB813    ;    //    sltiu x16 x23 -709      ====        sltiu a6, s7, -709
                                                  30'd    5096    : data = 32'h    01DE10B3    ;    //    sll x1 x28 x29      ====        sll ra, t3, t4
                                                  30'd    5097    : data = 32'h    4060D3B3    ;    //    sra x7 x1 x6      ====        sra t2, ra, t1
                                                  30'd    5098    : data = 32'h    0193D2B3    ;    //    srl x5 x7 x25      ====        srl t0, t2, s9
                                                  30'd    5099    : data = 32'h    00118D33    ;    //    add x26 x3 x1      ====        add s10, gp, ra
                                                  30'd    5100    : data = 32'h    D7398313    ;    //    addi x6 x19 -653      ====        addi t1, s3, -653
                                                  30'd    5101    : data = 32'h    09010A13    ;    //    addi x20 x2 144      ====        addi s4, sp, 144
                                                  30'd    5102    : data = 32'h    01426333    ;    //    or x6 x4 x20      ====        or t1, tp, s4
                                                  30'd    5103    : data = 32'h    40FFD6B3    ;    //    sra x13 x31 x15      ====        sra a3, t6, a5
                                                  30'd    5104    : data = 32'h    E93F4F93    ;    //    xori x31 x30 -365      ====        xori t6, t5, -365
                                                  30'd    5105    : data = 32'h    41F2DCB3    ;    //    sra x25 x5 x31      ====        sra s9, t0, t6
                                                  30'd    5106    : data = 32'h    009BAE33    ;    //    slt x28 x23 x9      ====        slt t3, s7, s1
                                                  30'd    5107    : data = 32'h    3BBAE313    ;    //    ori x6 x21 955      ====        ori t1, s5, 955
                                                  30'd    5108    : data = 32'h    01EA8433    ;    //    add x8 x21 x30      ====        add s0, s5, t5
                                                  30'd    5109    : data = 32'h    2FEDF993    ;    //    andi x19 x27 766      ====        andi s3, s11, 766
                                                  30'd    5110    : data = 32'h    1EDBA913    ;    //    slti x18 x23 493      ====        slti s2, s7, 493
                                                  30'd    5111    : data = 32'h    0198D593    ;    //    srli x11 x17 25      ====        srli a1, a7, 25
                                                  30'd    5112    : data = 32'h    C03BE413    ;    //    ori x8 x23 -1021      ====        ori s0, s7, -1021
                                                  30'd    5113    : data = 32'h    01BCC733    ;    //    xor x14 x25 x27      ====        xor a4, s9, s11
                                                  30'd    5114    : data = 32'h    00C32AB3    ;    //    slt x21 x6 x12      ====        slt s5, t1, a2
                                                  30'd    5115    : data = 32'h    00E21813    ;    //    slli x16 x4 14      ====        slli a6, tp, 14
                                                  30'd    5116    : data = 32'h    8F452293    ;    //    slti x5 x10 -1804      ====        slti t0, a0, -1804
                                                  30'd    5117    : data = 32'h    00E1C733    ;    //    xor x14 x3 x14      ====        xor a4, gp, a4
                                                  30'd    5118    : data = 32'h    22272097    ;    //    auipc x1 139890      ====        auipc ra, 139890
                                                  30'd    5119    : data = 32'h    00B794B3    ;    //    sll x9 x15 x11      ====        sll s1, a5, a1
                                                  30'd    5120    : data = 32'h    01095E93    ;    //    srli x29 x18 16      ====        srli t4, s2, 16
                                                  30'd    5121    : data = 32'h    01F9E433    ;    //    or x8 x19 x31      ====        or s0, s3, t6
                                                  30'd    5122    : data = 32'h    01E9BD33    ;    //    sltu x26 x19 x30      ====        sltu s10, s3, t5
                                                  30'd    5123    : data = 32'h    01CD5B33    ;    //    srl x22 x26 x28      ====        srl s6, s10, t3
                                                  30'd    5124    : data = 32'h    4020D033    ;    //    sra x0 x1 x2      ====        sra zero, ra, sp
                                                  30'd    5125    : data = 32'h    40FD5DB3    ;    //    sra x27 x26 x15      ====        sra s11, s10, a5
                                                  30'd    5126    : data = 32'h    0030FD33    ;    //    and x26 x1 x3      ====        and s10, ra, gp
                                                  30'd    5127    : data = 32'h    4129D693    ;    //    srai x13 x19 18      ====        srai a3, s3, 18
                                                  30'd    5128    : data = 32'h    40405333    ;    //    sra x6 x0 x4      ====        sra t1, zero, tp
                                                  30'd    5129    : data = 32'h    41DA8933    ;    //    sub x18 x21 x29      ====        sub s2, s5, t4
                                                  30'd    5130    : data = 32'h    40DB5093    ;    //    srai x1 x22 13      ====        srai ra, s6, 13
                                                  30'd    5131    : data = 32'h    00435713    ;    //    srli x14 x6 4      ====        srli a4, t1, 4
                                                  30'd    5132    : data = 32'h    413B5B33    ;    //    sra x22 x22 x19      ====        sra s6, s6, s3
                                                  30'd    5133    : data = 32'h    0A9D8793    ;    //    addi x15 x27 169      ====        addi a5, s11, 169
                                                  30'd    5134    : data = 32'h    EB420D13    ;    //    addi x26 x4 -332      ====        addi s10, tp, -332
                                                  30'd    5135    : data = 32'h    00791713    ;    //    slli x14 x18 7      ====        slli a4, s2, 7
                                                  30'd    5136    : data = 32'h    BE17E293    ;    //    ori x5 x15 -1055      ====        ori t0, a5, -1055
                                                  30'd    5137    : data = 32'h    5E358A93    ;    //    addi x21 x11 1507      ====        addi s5, a1, 1507
                                                  30'd    5138    : data = 32'h    407159B3    ;    //    sra x19 x2 x7      ====        sra s3, sp, t2
                                                  30'd    5139    : data = 32'h    01E71E33    ;    //    sll x28 x14 x30      ====        sll t3, a4, t5
                                                  30'd    5140    : data = 32'h    14748A93    ;    //    addi x21 x9 327      ====        addi s5, s1, 327
                                                  30'd    5141    : data = 32'h    00A93433    ;    //    sltu x8 x18 x10      ====        sltu s0, s2, a0
                                                  30'd    5142    : data = 32'h    5FC42393    ;    //    slti x7 x8 1532      ====        slti t2, s0, 1532
                                                  30'd    5143    : data = 32'h    004B9993    ;    //    slli x19 x23 4      ====        slli s3, s7, 4
                                                  30'd    5144    : data = 32'h    00E4D133    ;    //    srl x2 x9 x14      ====        srl sp, s1, a4
                                                  30'd    5145    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5146    : data = 32'h    7A6BEFB7    ;    //    lui x31 501438      ====        lui t6, 501438
                                                  30'd    5147    : data = 32'h    C4F9B913    ;    //    sltiu x18 x19 -945      ====        sltiu s2, s3, -945
                                                  30'd    5148    : data = 32'h    00FAED33    ;    //    or x26 x21 x15      ====        or s10, s5, a5
                                                  30'd    5149    : data = 32'h    C8ADAA13    ;    //    slti x20 x27 -886      ====        slti s4, s11, -886
                                                  30'd    5150    : data = 32'h    015CAD33    ;    //    slt x26 x25 x21      ====        slt s10, s9, s5
                                                  30'd    5151    : data = 32'h    008668B3    ;    //    or x17 x12 x8      ====        or a7, a2, s0
                                                  30'd    5152    : data = 32'h    7383FE13    ;    //    andi x28 x7 1848      ====        andi t3, t2, 1848
                                                  30'd    5153    : data = 32'h    40765033    ;    //    sra x0 x12 x7      ====        sra zero, a2, t2
                                                  30'd    5154    : data = 32'h    00375593    ;    //    srli x11 x14 3      ====        srli a1, a4, 3
                                                  30'd    5155    : data = 32'h    00827BB3    ;    //    and x23 x4 x8      ====        and s7, tp, s0
                                                  30'd    5156    : data = 32'h    011A74B3    ;    //    and x9 x20 x17      ====        and s1, s4, a7
                                                  30'd    5157    : data = 32'h    F00FF1B7    ;    //    lui x3 983295      ====        lui gp, 983295
                                                  30'd    5158    : data = 32'h    403402B3    ;    //    sub x5 x8 x3      ====        sub t0, s0, gp
                                                  30'd    5159    : data = 32'h    014BF1B3    ;    //    and x3 x23 x20      ====        and gp, s7, s4
                                                  30'd    5160    : data = 32'h    410AD313    ;    //    srai x6 x21 16      ====        srai t1, s5, 16
                                                  30'd    5161    : data = 32'h    01031813    ;    //    slli x16 x6 16      ====        slli a6, t1, 16
                                                  30'd    5162    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5163    : data = 32'h    641E2113    ;    //    slti x2 x28 1601      ====        slti sp, t3, 1601
                                                  30'd    5164    : data = 32'h    8DE7CC13    ;    //    xori x24 x15 -1826      ====        xori s8, a5, -1826
                                                  30'd    5165    : data = 32'h    003D1333    ;    //    sll x6 x26 x3      ====        sll t1, s10, gp
                                                  30'd    5166    : data = 32'h    0B250393    ;    //    addi x7 x10 178      ====        addi t2, a0, 178
                                                  30'd    5167    : data = 32'h    002E5B33    ;    //    srl x22 x28 x2      ====        srl s6, t3, sp
                                                  30'd    5168    : data = 32'h    3A08E113    ;    //    ori x2 x17 928      ====        ori sp, a7, 928
                                                  30'd    5169    : data = 32'h    C4E72493    ;    //    slti x9 x14 -946      ====        slti s1, a4, -946
                                                  30'd    5170    : data = 32'h    0178DCB3    ;    //    srl x25 x17 x23      ====        srl s9, a7, s7
                                                  30'd    5171    : data = 32'h    4006D633    ;    //    sra x12 x13 x0      ====        sra a2, a3, zero
                                                  30'd    5172    : data = 32'h    41D95113    ;    //    srai x2 x18 29      ====        srai sp, s2, 29
                                                  30'd    5173    : data = 32'h    01C69613    ;    //    slli x12 x13 28      ====        slli a2, a3, 28
                                                  30'd    5174    : data = 32'h    401E5013    ;    //    srai x0 x28 1      ====        srai zero, t3, 1
                                                  30'd    5175    : data = 32'h    2D1FF113    ;    //    andi x2 x31 721      ====        andi sp, t6, 721
                                                  30'd    5176    : data = 32'h    40CED813    ;    //    srai x16 x29 12      ====        srai a6, t4, 12
                                                  30'd    5177    : data = 32'h    417BDCB3    ;    //    sra x25 x23 x23      ====        sra s9, s7, s7
                                                  30'd    5178    : data = 32'h    01A93033    ;    //    sltu x0 x18 x26      ====        sltu zero, s2, s10
                                                  30'd    5179    : data = 32'h    0032EEB3    ;    //    or x29 x5 x3      ====        or t4, t0, gp
                                                  30'd    5180    : data = 32'h    65CC4113    ;    //    xori x2 x24 1628      ====        xori sp, s8, 1628
                                                  30'd    5181    : data = 32'h    0107D733    ;    //    srl x14 x15 x16      ====        srl a4, a5, a6
                                                  30'd    5182    : data = 32'h    0158C033    ;    //    xor x0 x17 x21      ====        xor zero, a7, s5
                                                  30'd    5183    : data = 32'h    01907A33    ;    //    and x20 x0 x25      ====        and s4, zero, s9
                                                  30'd    5184    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5185    : data = 32'h    41118433    ;    //    sub x8 x3 x17      ====        sub s0, gp, a7
                                                  30'd    5186    : data = 32'h    019C44B3    ;    //    xor x9 x24 x25      ====        xor s1, s8, s9
                                                  30'd    5187    : data = 32'h    4D04C093    ;    //    xori x1 x9 1232      ====        xori ra, s1, 1232
                                                  30'd    5188    : data = 32'h    14407B17    ;    //    auipc x22 82951      ====        auipc s6, 82951
                                                  30'd    5189    : data = 32'h    01039313    ;    //    slli x6 x7 16      ====        slli t1, t2, 16
                                                  30'd    5190    : data = 32'h    018A18B3    ;    //    sll x17 x20 x24      ====        sll a7, s4, s8
                                                  30'd    5191    : data = 32'h    8DBE0117    ;    //    auipc x2 580576      ====        auipc sp, 580576
                                                  30'd    5192    : data = 32'h    41D55D93    ;    //    srai x27 x10 29      ====        srai s11, a0, 29
                                                  30'd    5193    : data = 32'h    10E08A93    ;    //    addi x21 x1 270      ====        addi s5, ra, 270
                                                  30'd    5194    : data = 32'h    5B768013    ;    //    addi x0 x13 1463      ====        addi zero, a3, 1463
                                                  30'd    5195    : data = 32'h    01ED5733    ;    //    srl x14 x26 x30      ====        srl a4, s10, t5
                                                  30'd    5196    : data = 32'h    B753ED13    ;    //    ori x26 x7 -1163      ====        ori s10, t2, -1163
                                                  30'd    5197    : data = 32'h    F22F0613    ;    //    addi x12 x30 -222      ====        addi a2, t5, -222
                                                  30'd    5198    : data = 32'h    996A8793    ;    //    addi x15 x21 -1642      ====        addi a5, s5, -1642
                                                  30'd    5199    : data = 32'h    00CC0FB3    ;    //    add x31 x24 x12      ====        add t6, s8, a2
                                                  30'd    5200    : data = 32'h    58A67B13    ;    //    andi x22 x12 1418      ====        andi s6, a2, 1418
                                                  30'd    5201    : data = 32'h    40A80C33    ;    //    sub x24 x16 x10      ====        sub s8, a6, a0
                                                  30'd    5202    : data = 32'h    00EA9EB3    ;    //    sll x29 x21 x14      ====        sll t4, s5, a4
                                                  30'd    5203    : data = 32'h    1A2C6197    ;    //    auipc x3 107206      ====        auipc gp, 107206
                                                  30'd    5204    : data = 32'h    416F0C33    ;    //    sub x24 x30 x22      ====        sub s8, t5, s6
                                                  30'd    5205    : data = 32'h    000D5893    ;    //    srli x17 x26 0      ====        srli a7, s10, 0
                                                  30'd    5206    : data = 32'h    40C05B13    ;    //    srai x22 x0 12      ====        srai s6, zero, 12
                                                  30'd    5207    : data = 32'h    40878033    ;    //    sub x0 x15 x8      ====        sub zero, a5, s0
                                                  30'd    5208    : data = 32'h    00068A33    ;    //    add x20 x13 x0      ====        add s4, a3, zero
                                                  30'd    5209    : data = 32'h    40638033    ;    //    sub x0 x7 x6      ====        sub zero, t2, t1
                                                  30'd    5210    : data = 32'h    C3212793    ;    //    slti x15 x2 -974      ====        slti a5, sp, -974
                                                  30'd    5211    : data = 32'h    013468B3    ;    //    or x17 x8 x19      ====        or a7, s0, s3
                                                  30'd    5212    : data = 32'h    41B1D4B3    ;    //    sra x9 x3 x27      ====        sra s1, gp, s11
                                                  30'd    5213    : data = 32'h    B0B644B7    ;    //    lui x9 723812      ====        lui s1, 723812
                                                  30'd    5214    : data = 32'h    016D0E33    ;    //    add x28 x26 x22      ====        add t3, s10, s6
                                                  30'd    5215    : data = 32'h    010F50B3    ;    //    srl x1 x30 x16      ====        srl ra, t5, a6
                                                  30'd    5216    : data = 32'h    A9762F93    ;    //    slti x31 x12 -1385      ====        slti t6, a2, -1385
                                                  30'd    5217    : data = 32'h    471E6E13    ;    //    ori x28 x28 1137      ====        ori t3, t3, 1137
                                                  30'd    5218    : data = 32'h    40D98D33    ;    //    sub x26 x19 x13      ====        sub s10, s3, a3
                                                  30'd    5219    : data = 32'h    3A9EA493    ;    //    slti x9 x29 937      ====        slti s1, t4, 937
                                                  30'd    5220    : data = 32'h    018D21B3    ;    //    slt x3 x26 x24      ====        slt gp, s10, s8
                                                  30'd    5221    : data = 32'h    01A94B33    ;    //    xor x22 x18 x26      ====        xor s6, s2, s10
                                                  30'd    5222    : data = 32'h    00D94FB3    ;    //    xor x31 x18 x13      ====        xor t6, s2, a3
                                                  30'd    5223    : data = 32'h    011BFCB3    ;    //    and x25 x23 x17      ====        and s9, s7, a7
                                                  30'd    5224    : data = 32'h    41FB86B3    ;    //    sub x13 x23 x31      ====        sub a3, s7, t6
                                                  30'd    5225    : data = 32'h    00A2A8B3    ;    //    slt x17 x5 x10      ====        slt a7, t0, a0
                                                  30'd    5226    : data = 32'h    01001B93    ;    //    slli x23 x0 16      ====        slli s7, zero, 16
                                                  30'd    5227    : data = 32'h    2BDA0D13    ;    //    addi x26 x20 701      ====        addi s10, s4, 701
                                                  30'd    5228    : data = 32'h    406E8EB3    ;    //    sub x29 x29 x6      ====        sub t4, t4, t1
                                                  30'd    5229    : data = 32'h    00807AB3    ;    //    and x21 x0 x8      ====        and s5, zero, s0
                                                  30'd    5230    : data = 32'h    1C9E7013    ;    //    andi x0 x28 457      ====        andi zero, t3, 457
                                                  30'd    5231    : data = 32'h    41158333    ;    //    sub x6 x11 x17      ====        sub t1, a1, a7
                                                  30'd    5232    : data = 32'h    401B52B3    ;    //    sra x5 x22 x1      ====        sra t0, s6, ra
                                                  30'd    5233    : data = 32'h    74D139B7    ;    //    lui x19 478483      ====        lui s3, 478483
                                                  30'd    5234    : data = 32'h    E4628337    ;    //    lui x6 935464      ====        lui t1, 935464
                                                  30'd    5235    : data = 32'h    B8EA47B7    ;    //    lui x15 757412      ====        lui a5, 757412
                                                  30'd    5236    : data = 32'h    0088D293    ;    //    srli x5 x17 8      ====        srli t0, a7, 8
                                                  30'd    5237    : data = 32'h    C5FE3013    ;    //    sltiu x0 x28 -929      ====        sltiu zero, t3, -929
                                                  30'd    5238    : data = 32'h    0193CAB3    ;    //    xor x21 x7 x25      ====        xor s5, t2, s9
                                                  30'd    5239    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5240    : data = 32'h    0092D793    ;    //    srli x15 x5 9      ====        srli a5, t0, 9
                                                  30'd    5241    : data = 32'h    66227613    ;    //    andi x12 x4 1634      ====        andi a2, tp, 1634
                                                  30'd    5242    : data = 32'h    01B49733    ;    //    sll x14 x9 x27      ====        sll a4, s1, s11
                                                  30'd    5243    : data = 32'h    696C2A13    ;    //    slti x20 x24 1686      ====        slti s4, s8, 1686
                                                  30'd    5244    : data = 32'h    2101A793    ;    //    slti x15 x3 528      ====        slti a5, gp, 528
                                                  30'd    5245    : data = 32'h    7CEC4193    ;    //    xori x3 x24 1998      ====        xori gp, s8, 1998
                                                  30'd    5246    : data = 32'h    40F302B3    ;    //    sub x5 x6 x15      ====        sub t0, t1, a5
                                                  30'd    5247    : data = 32'h    41635793    ;    //    srai x15 x6 22      ====        srai a5, t1, 22
                                                  30'd    5248    : data = 32'h    005D2CB3    ;    //    slt x25 x26 x5      ====        slt s9, s10, t0
                                                  30'd    5249    : data = 32'h    0133DF93    ;    //    srli x31 x7 19      ====        srli t6, t2, 19
                                                  30'd    5250    : data = 32'h    0020E333    ;    //    or x6 x1 x2      ====        or t1, ra, sp
                                                  30'd    5251    : data = 32'h    5F0B2B17    ;    //    auipc x22 389298      ====        auipc s6, 389298
                                                  30'd    5252    : data = 32'h    0089D013    ;    //    srli x0 x19 8      ====        srli zero, s3, 8
                                                  30'd    5253    : data = 32'h    415DD413    ;    //    srai x8 x27 21      ====        srai s0, s11, 21
                                                  30'd    5254    : data = 32'h    413CD333    ;    //    sra x6 x25 x19      ====        sra t1, s9, s3
                                                  30'd    5255    : data = 32'h    00A66433    ;    //    or x8 x12 x10      ====        or s0, a2, a0
                                                  30'd    5256    : data = 32'h    003EDE33    ;    //    srl x28 x29 x3      ====        srl t3, t4, gp
                                                  30'd    5257    : data = 32'h    B8F6F113    ;    //    andi x2 x13 -1137      ====        andi sp, a3, -1137
                                                  30'd    5258    : data = 32'h    00CE9DB3    ;    //    sll x27 x29 x12      ====        sll s11, t4, a2
                                                  30'd    5259    : data = 32'h    781B7E13    ;    //    andi x28 x22 1921      ====        andi t3, s6, 1921
                                                  30'd    5260    : data = 32'h    411B85B3    ;    //    sub x11 x23 x17      ====        sub a1, s7, a7
                                                  30'd    5261    : data = 32'h    00AA5B13    ;    //    srli x22 x20 10      ====        srli s6, s4, 10
                                                  30'd    5262    : data = 32'h    012496B3    ;    //    sll x13 x9 x18      ====        sll a3, s1, s2
                                                  30'd    5263    : data = 32'h    41965713    ;    //    srai x14 x12 25      ====        srai a4, a2, 25
                                                  30'd    5264    : data = 32'h    01A6D733    ;    //    srl x14 x13 x26      ====        srl a4, a3, s10
                                                  30'd    5265    : data = 32'h    12AB4713    ;    //    xori x14 x22 298      ====        xori a4, s6, 298
                                                  30'd    5266    : data = 32'h    01507D33    ;    //    and x26 x0 x21      ====        and s10, zero, s5
                                                  30'd    5267    : data = 32'h    4A874DB7    ;    //    lui x27 305268      ====        lui s11, 305268
                                                  30'd    5268    : data = 32'h    01EEB6B3    ;    //    sltu x13 x29 x30      ====        sltu a3, t4, t5
                                                  30'd    5269    : data = 32'h    008670B3    ;    //    and x1 x12 x8      ====        and ra, a2, s0
                                                  30'd    5270    : data = 32'h    00DE7CB3    ;    //    and x25 x28 x13      ====        and s9, t3, a3
                                                  30'd    5271    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5272    : data = 32'h    05286C13    ;    //    ori x24 x16 82      ====        ori s8, a6, 82
                                                  30'd    5273    : data = 32'h    0038A833    ;    //    slt x16 x17 x3      ====        slt a6, a7, gp
                                                  30'd    5274    : data = 32'h    88F66F93    ;    //    ori x31 x12 -1905      ====        ori t6, a2, -1905
                                                  30'd    5275    : data = 32'h    17F7AA93    ;    //    slti x21 x15 383      ====        slti s5, a5, 383
                                                  30'd    5276    : data = 32'h    22E2DDB7    ;    //    lui x27 142893      ====        lui s11, 142893
                                                  30'd    5277    : data = 32'h    BB618C93    ;    //    addi x25 x3 -1098      ====        addi s9, gp, -1098
                                                  30'd    5278    : data = 32'h    01F47A33    ;    //    and x20 x8 x31      ====        and s4, s0, t6
                                                  30'd    5279    : data = 32'h    80E4E313    ;    //    ori x6 x9 -2034      ====        ori t1, s1, -2034
                                                  30'd    5280    : data = 32'h    41518B33    ;    //    sub x22 x3 x21      ====        sub s6, gp, s5
                                                  30'd    5281    : data = 32'h    007A03B3    ;    //    add x7 x20 x7      ====        add t2, s4, t2
                                                  30'd    5282    : data = 32'h    0017B433    ;    //    sltu x8 x15 x1      ====        sltu s0, a5, ra
                                                  30'd    5283    : data = 32'h    7BADDFB7    ;    //    lui x31 506589      ====        lui t6, 506589
                                                  30'd    5284    : data = 32'h    04CE2413    ;    //    slti x8 x28 76      ====        slti s0, t3, 76
                                                  30'd    5285    : data = 32'h    41FC8CB3    ;    //    sub x25 x25 x31      ====        sub s9, s9, t6
                                                  30'd    5286    : data = 32'h    007BDF93    ;    //    srli x31 x23 7      ====        srli t6, s7, 7
                                                  30'd    5287    : data = 32'h    406706B3    ;    //    sub x13 x14 x6      ====        sub a3, a4, t1
                                                  30'd    5288    : data = 32'h    005C1433    ;    //    sll x8 x24 x5      ====        sll s0, s8, t0
                                                  30'd    5289    : data = 32'h    1D092197    ;    //    auipc x3 118930      ====        auipc gp, 118930
                                                  30'd    5290    : data = 32'h    012C33B3    ;    //    sltu x7 x24 x18      ====        sltu t2, s8, s2
                                                  30'd    5291    : data = 32'h    01AB3BB3    ;    //    sltu x23 x22 x26      ====        sltu s7, s6, s10
                                                  30'd    5292    : data = 32'h    F762B993    ;    //    sltiu x19 x5 -138      ====        sltiu s3, t0, -138
                                                  30'd    5293    : data = 32'h    009E2EB3    ;    //    slt x29 x28 x9      ====        slt t4, t3, s1
                                                  30'd    5294    : data = 32'h    414A8833    ;    //    sub x16 x21 x20      ====        sub a6, s5, s4
                                                  30'd    5295    : data = 32'h    B7DE6917    ;    //    auipc x18 753126      ====        auipc s2, 753126
                                                  30'd    5296    : data = 32'h    DBA4C013    ;    //    xori x0 x9 -582      ====        xori zero, s1, -582
                                                  30'd    5297    : data = 32'h    16A33413    ;    //    sltiu x8 x6 362      ====        sltiu s0, t1, 362
                                                  30'd    5298    : data = 32'h    011FFCB3    ;    //    and x25 x31 x17      ====        and s9, t6, a7
                                                  30'd    5299    : data = 32'h    C7502193    ;    //    slti x3 x0 -907      ====        slti gp, zero, -907
                                                  30'd    5300    : data = 32'h    3FEBAA13    ;    //    slti x20 x23 1022      ====        slti s4, s7, 1022
                                                  30'd    5301    : data = 32'h    01AF8A33    ;    //    add x20 x31 x26      ====        add s4, t6, s10
                                                  30'd    5302    : data = 32'h    016F0EB3    ;    //    add x29 x30 x22      ====        add t4, t5, s6
                                                  30'd    5303    : data = 32'h    00D46AB3    ;    //    or x21 x8 x13      ====        or s5, s0, a3
                                                  30'd    5304    : data = 32'h    5D2BC813    ;    //    xori x16 x23 1490      ====        xori a6, s7, 1490
                                                  30'd    5305    : data = 32'h    41395633    ;    //    sra x12 x18 x19      ====        sra a2, s2, s3
                                                  30'd    5306    : data = 32'h    01838B33    ;    //    add x22 x7 x24      ====        add s6, t2, s8
                                                  30'd    5307    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5308    : data = 32'h    017A40B3    ;    //    xor x1 x20 x23      ====        xor ra, s4, s7
                                                  30'd    5309    : data = 32'h    10BAAB37    ;    //    lui x22 68522      ====        lui s6, 68522
                                                  30'd    5310    : data = 32'h    003E16B3    ;    //    sll x13 x28 x3      ====        sll a3, t3, gp
                                                  30'd    5311    : data = 32'h    01C22D33    ;    //    slt x26 x4 x28      ====        slt s10, tp, t3
                                                  30'd    5312    : data = 32'h    41A20E33    ;    //    sub x28 x4 x26      ====        sub t3, tp, s10
                                                  30'd    5313    : data = 32'h    A4017293    ;    //    andi x5 x2 -1472      ====        andi t0, sp, -1472
                                                  30'd    5314    : data = 32'h    40C080B3    ;    //    sub x1 x1 x12      ====        sub ra, ra, a2
                                                  30'd    5315    : data = 32'h    01FCD193    ;    //    srli x3 x25 31      ====        srli gp, s9, 31
                                                  30'd    5316    : data = 32'h    00243E33    ;    //    sltu x28 x8 x2      ====        sltu t3, s0, sp
                                                  30'd    5317    : data = 32'h    0845CA13    ;    //    xori x20 x11 132      ====        xori s4, a1, 132
                                                  30'd    5318    : data = 32'h    EC52EC93    ;    //    ori x25 x5 -315      ====        ori s9, t0, -315
                                                  30'd    5319    : data = 32'h    01E7E4B3    ;    //    or x9 x15 x30      ====        or s1, a5, t5
                                                  30'd    5320    : data = 32'h    825CB793    ;    //    sltiu x15 x25 -2011      ====        sltiu a5, s9, -2011
                                                  30'd    5321    : data = 32'h    412502B3    ;    //    sub x5 x10 x18      ====        sub t0, a0, s2
                                                  30'd    5322    : data = 32'h    41975313    ;    //    srai x6 x14 25      ====        srai t1, a4, 25
                                                  30'd    5323    : data = 32'h    01E2DCB3    ;    //    srl x25 x5 x30      ====        srl s9, t0, t5
                                                  30'd    5324    : data = 32'h    00D1D893    ;    //    srli x17 x3 13      ====        srli a7, gp, 13
                                                  30'd    5325    : data = 32'h    00695B13    ;    //    srli x22 x18 6      ====        srli s6, s2, 6
                                                  30'd    5326    : data = 32'h    00A9ABB3    ;    //    slt x23 x19 x10      ====        slt s7, s3, a0
                                                  30'd    5327    : data = 32'h    008CDB33    ;    //    srl x22 x25 x8      ====        srl s6, s9, s0
                                                  30'd    5328    : data = 32'h    0064E6B3    ;    //    or x13 x9 x6      ====        or a3, s1, t1
                                                  30'd    5329    : data = 32'h    01392FB3    ;    //    slt x31 x18 x19      ====        slt t6, s2, s3
                                                  30'd    5330    : data = 32'h    6D9479B7    ;    //    lui x19 448839      ====        lui s3, 448839
                                                  30'd    5331    : data = 32'h    0082AFB3    ;    //    slt x31 x5 x8      ====        slt t6, t0, s0
                                                  30'd    5332    : data = 32'h    0123E033    ;    //    or x0 x7 x18      ====        or zero, t2, s2
                                                  30'd    5333    : data = 32'h    00369933    ;    //    sll x18 x13 x3      ====        sll s2, a3, gp
                                                  30'd    5334    : data = 32'h    01B13CB3    ;    //    sltu x25 x2 x27      ====        sltu s9, sp, s11
                                                  30'd    5335    : data = 32'h    41B85893    ;    //    srai x17 x16 27      ====        srai a7, a6, 27
                                                  30'd    5336    : data = 32'h    01809933    ;    //    sll x18 x1 x24      ====        sll s2, ra, s8
                                                  30'd    5337    : data = 32'h    40AED413    ;    //    srai x8 x29 10      ====        srai s0, t4, 10
                                                  30'd    5338    : data = 32'h    40B3D813    ;    //    srai x16 x7 11      ====        srai a6, t2, 11
                                                  30'd    5339    : data = 32'h    7B286E17    ;    //    auipc x28 504454      ====        auipc t3, 504454
                                                  30'd    5340    : data = 32'h    010AD9B3    ;    //    srl x19 x21 x16      ====        srl s3, s5, a6
                                                  30'd    5341    : data = 32'h    EE076693    ;    //    ori x13 x14 -288      ====        ori a3, a4, -288
                                                  30'd    5342    : data = 32'h    00492A33    ;    //    slt x20 x18 x4      ====        slt s4, s2, tp
                                                  30'd    5343    : data = 32'h    41520D33    ;    //    sub x26 x4 x21      ====        sub s10, tp, s5
                                                  30'd    5344    : data = 32'h    01121733    ;    //    sll x14 x4 x17      ====        sll a4, tp, a7
                                                  30'd    5345    : data = 32'h    F6D92913    ;    //    slti x18 x18 -147      ====        slti s2, s2, -147
                                                  30'd    5346    : data = 32'h    01E884B3    ;    //    add x9 x17 x30      ====        add s1, a7, t5
                                                  30'd    5347    : data = 32'h    25F14993    ;    //    xori x19 x2 607      ====        xori s3, sp, 607
                                                  30'd    5348    : data = 32'h    2E146B93    ;    //    ori x23 x8 737      ====        ori s7, s0, 737
                                                  30'd    5349    : data = 32'h    3B52E593    ;    //    ori x11 x5 949      ====        ori a1, t0, 949
                                                  30'd    5350    : data = 32'h    018381B3    ;    //    add x3 x7 x24      ====        add gp, t2, s8
                                                  30'd    5351    : data = 32'h    003E1E33    ;    //    sll x28 x28 x3      ====        sll t3, t3, gp
                                                  30'd    5352    : data = 32'h    7FD92A13    ;    //    slti x20 x18 2045      ====        slti s4, s2, 2045
                                                  30'd    5353    : data = 32'h    D028CCB7    ;    //    lui x25 852620      ====        lui s9, 852620
                                                  30'd    5354    : data = 32'h    999C4793    ;    //    xori x15 x24 -1639      ====        xori a5, s8, -1639
                                                  30'd    5355    : data = 32'h    4069DB13    ;    //    srai x22 x19 6      ====        srai s6, s3, 6
                                                  30'd    5356    : data = 32'h    D0120913    ;    //    addi x18 x4 -767      ====        addi s2, tp, -767
                                                  30'd    5357    : data = 32'h    00C75D93    ;    //    srli x27 x14 12      ====        srli s11, a4, 12
                                                  30'd    5358    : data = 32'h    41CA84B3    ;    //    sub x9 x21 x28      ====        sub s1, s5, t3
                                                  30'd    5359    : data = 32'h    E8683113    ;    //    sltiu x2 x16 -378      ====        sltiu sp, a6, -378
                                                  30'd    5360    : data = 32'h    0208A717    ;    //    auipc x14 8330      ====        auipc a4, 8330
                                                  30'd    5361    : data = 32'h    4AC3F013    ;    //    andi x0 x7 1196      ====        andi zero, t2, 1196
                                                  30'd    5362    : data = 32'h    010B5033    ;    //    srl x0 x22 x16      ====        srl zero, s6, a6
                                                  30'd    5363    : data = 32'h    001E68B3    ;    //    or x17 x28 x1      ====        or a7, t3, ra
                                                  30'd    5364    : data = 32'h    41440B33    ;    //    sub x22 x8 x20      ====        sub s6, s0, s4
                                                  30'd    5365    : data = 32'h    EBC3CA13    ;    //    xori x20 x7 -324      ====        xori s4, t2, -324
                                                  30'd    5366    : data = 32'h    000962B3    ;    //    or x5 x18 x0      ====        or t0, s2, zero
                                                  30'd    5367    : data = 32'h    414BD293    ;    //    srai x5 x23 20      ====        srai t0, s7, 20
                                                  30'd    5368    : data = 32'h    40660033    ;    //    sub x0 x12 x6      ====        sub zero, a2, t1
                                                  30'd    5369    : data = 32'h    01FBA3B3    ;    //    slt x7 x23 x31      ====        slt t2, s7, t6
                                                  30'd    5370    : data = 32'h    B0A4F613    ;    //    andi x12 x9 -1270      ====        andi a2, s1, -1270
                                                  30'd    5371    : data = 32'h    5A7FA313    ;    //    slti x6 x31 1447      ====        slti t1, t6, 1447
                                                  30'd    5372    : data = 32'h    0072BB33    ;    //    sltu x22 x5 x7      ====        sltu s6, t0, t2
                                                  30'd    5373    : data = 32'h    01F6F5B3    ;    //    and x11 x13 x31      ====        and a1, a3, t6
                                                  30'd    5374    : data = 32'h    00DE1633    ;    //    sll x12 x28 x13      ====        sll a2, t3, a3
                                                  30'd    5375    : data = 32'h    01D9E6B3    ;    //    or x13 x19 x29      ====        or a3, s3, t4
                                                  30'd    5376    : data = 32'h    401DD013    ;    //    srai x0 x27 1      ====        srai zero, s11, 1
                                                  30'd    5377    : data = 32'h    AD869A97    ;    //    auipc x21 710761      ====        auipc s5, 710761
                                                  30'd    5378    : data = 32'h    01BC1593    ;    //    slli x11 x24 27      ====        slli a1, s8, 27
                                                  30'd    5379    : data = 32'h    0086BDB3    ;    //    sltu x27 x13 x8      ====        sltu s11, a3, s0
                                                  30'd    5380    : data = 32'h    41180133    ;    //    sub x2 x16 x17      ====        sub sp, a6, a7
                                                  30'd    5381    : data = 32'h    C3BCCDB7    ;    //    lui x27 801740      ====        lui s11, 801740
                                                  30'd    5382    : data = 32'h    0DC58B93    ;    //    addi x23 x11 220      ====        addi s7, a1, 220
                                                  30'd    5383    : data = 32'h    D57DFF93    ;    //    andi x31 x27 -681      ====        andi t6, s11, -681
                                                  30'd    5384    : data = 32'h    015BD4B3    ;    //    srl x9 x23 x21      ====        srl s1, s7, s5
                                                  30'd    5385    : data = 32'h    002C66B3    ;    //    or x13 x24 x2      ====        or a3, s8, sp
                                                  30'd    5386    : data = 32'h    01C87033    ;    //    and x0 x16 x28      ====        and zero, a6, t3
                                                  30'd    5387    : data = 32'h    26F4BC37    ;    //    lui x24 159563      ====        lui s8, 159563
                                                  30'd    5388    : data = 32'h    5ED25797    ;    //    auipc x15 388389      ====        auipc a5, 388389
                                                  30'd    5389    : data = 32'h    10CCEC13    ;    //    ori x24 x25 268      ====        ori s8, s9, 268
                                                  30'd    5390    : data = 32'h    00A178B3    ;    //    and x17 x2 x10      ====        and a7, sp, a0
                                                  30'd    5391    : data = 32'h    00BA4833    ;    //    xor x16 x20 x11      ====        xor a6, s4, a1
                                                  30'd    5392    : data = 32'h    9F30FD17    ;    //    auipc x26 652047      ====        auipc s10, 652047
                                                  30'd    5393    : data = 32'h    E5190393    ;    //    addi x7 x18 -431      ====        addi t2, s2, -431
                                                  30'd    5394    : data = 32'h    01A180B3    ;    //    add x1 x3 x26      ====        add ra, gp, s10
                                                  30'd    5395    : data = 32'h    017DA0B3    ;    //    slt x1 x27 x23      ====        slt ra, s11, s7
                                                  30'd    5396    : data = 32'h    939BB097    ;    //    auipc x1 604603      ====        auipc ra, 604603
                                                  30'd    5397    : data = 32'h    58D53013    ;    //    sltiu x0 x10 1421      ====        sltiu zero, a0, 1421
                                                  30'd    5398    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5399    : data = 32'h    00702BB3    ;    //    slt x23 x0 x7      ====        slt s7, zero, t2
                                                  30'd    5400    : data = 32'h    27FDBE97    ;    //    auipc x29 163803      ====        auipc t4, 163803
                                                  30'd    5401    : data = 32'h    01B77833    ;    //    and x16 x14 x27      ====        and a6, a4, s11
                                                  30'd    5402    : data = 32'h    40B50D33    ;    //    sub x26 x10 x11      ====        sub s10, a0, a1
                                                  30'd    5403    : data = 32'h    003F1D33    ;    //    sll x26 x30 x3      ====        sll s10, t5, gp
                                                  30'd    5404    : data = 32'h    0158DDB3    ;    //    srl x27 x17 x21      ====        srl s11, a7, s5
                                                  30'd    5405    : data = 32'h    013EDDB3    ;    //    srl x27 x29 x19      ====        srl s11, t4, s3
                                                  30'd    5406    : data = 32'h    EBA84C13    ;    //    xori x24 x16 -326      ====        xori s8, a6, -326
                                                  30'd    5407    : data = 32'h    400D54B3    ;    //    sra x9 x26 x0      ====        sra s1, s10, zero
                                                  30'd    5408    : data = 32'h    00045733    ;    //    srl x14 x8 x0      ====        srl a4, s0, zero
                                                  30'd    5409    : data = 32'h    0047CE33    ;    //    xor x28 x15 x4      ====        xor t3, a5, tp
                                                  30'd    5410    : data = 32'h    9B4134B7    ;    //    lui x9 635923      ====        lui s1, 635923
                                                  30'd    5411    : data = 32'h    0122F133    ;    //    and x2 x5 x18      ====        and sp, t0, s2
                                                  30'd    5412    : data = 32'h    011F2133    ;    //    slt x2 x30 x17      ====        slt sp, t5, a7
                                                  30'd    5413    : data = 32'h    87DAA313    ;    //    slti x6 x21 -1923      ====        slti t1, s5, -1923
                                                  30'd    5414    : data = 32'h    CEB2FB97    ;    //    auipc x23 846639      ====        auipc s7, 846639
                                                  30'd    5415    : data = 32'h    01A5B9B3    ;    //    sltu x19 x11 x26      ====        sltu s3, a1, s10
                                                  30'd    5416    : data = 32'h    013F35B3    ;    //    sltu x11 x30 x19      ====        sltu a1, t5, s3
                                                  30'd    5417    : data = 32'h    6E76C713    ;    //    xori x14 x13 1767      ====        xori a4, a3, 1767
                                                  30'd    5418    : data = 32'h    329BED93    ;    //    ori x27 x23 809      ====        ori s11, s7, 809
                                                  30'd    5419    : data = 32'h    00CEDBB3    ;    //    srl x23 x29 x12      ====        srl s7, t4, a2
                                                  30'd    5420    : data = 32'h    38A88413    ;    //    addi x8 x17 906      ====        addi s0, a7, 906
                                                  30'd    5421    : data = 32'h    873A97B7    ;    //    lui x15 553897      ====        lui a5, 553897
                                                  30'd    5422    : data = 32'h    418B5A13    ;    //    srai x20 x22 24      ====        srai s4, s6, 24
                                                  30'd    5423    : data = 32'h    01293A33    ;    //    sltu x20 x18 x18      ====        sltu s4, s2, s2
                                                  30'd    5424    : data = 32'h    00CE1F93    ;    //    slli x31 x28 12      ====        slli t6, t3, 12
                                                  30'd    5425    : data = 32'h    00AB05B3    ;    //    add x11 x22 x10      ====        add a1, s6, a0
                                                  30'd    5426    : data = 32'h    01BB61B3    ;    //    or x3 x22 x27      ====        or gp, s6, s11
                                                  30'd    5427    : data = 32'h    41978B33    ;    //    sub x22 x15 x25      ====        sub s6, a5, s9
                                                  30'd    5428    : data = 32'h    00939B13    ;    //    slli x22 x7 9      ====        slli s6, t2, 9
                                                  30'd    5429    : data = 32'h    3177B313    ;    //    sltiu x6 x15 791      ====        sltiu t1, a5, 791
                                                  30'd    5430    : data = 32'h    00A02933    ;    //    slt x18 x0 x10      ====        slt s2, zero, a0
                                                  30'd    5431    : data = 32'h    006F5E33    ;    //    srl x28 x30 x6      ====        srl t3, t5, t1
                                                  30'd    5432    : data = 32'h    FFF00413    ;    //    addi x8 x0 -1      ====        li s0, 0xffffffff #start riscv_int_numeric_corner_stream_31
                                                  30'd    5433    : data = 32'h    00000A93    ;    //    addi x21 x0 0      ====        li s5, 0x0
                                                  30'd    5434    : data = 32'h    5ECDCDB7    ;    //    lui x27 388316      ====        li s11, 0x5ecdc4b7
                                                  30'd    5435    : data = 32'h    4B7D8D93    ;    //    addi x27 x27 1207      ====        li s11, 0x5ecdc4b7
                                                  30'd    5436    : data = 32'h    00000713    ;    //    addi x14 x0 0      ====        li a4, 0x0
                                                  30'd    5437    : data = 32'h    FFF00893    ;    //    addi x17 x0 -1      ====        li a7, 0xffffffff
                                                  30'd    5438    : data = 32'h    DDEF91B7    ;    //    lui x3 909049      ====        li gp, 0xddef9163
                                                  30'd    5439    : data = 32'h    16318193    ;    //    addi x3 x3 355      ====        li gp, 0xddef9163
                                                  30'd    5440    : data = 32'h    80000A37    ;    //    lui x20 524288      ====        li s4, 0x80000000
                                                  30'd    5441    : data = 32'h    000A0A13    ;    //    addi x20 x20 0      ====        li s4, 0x80000000
                                                  30'd    5442    : data = 32'h    9C18F137    ;    //    lui x2 639375      ====        li sp, 0x9c18ef92
                                                  30'd    5443    : data = 32'h    F9210113    ;    //    addi x2 x2 -110      ====        li sp, 0x9c18ef92
                                                  30'd    5444    : data = 32'h    5BE2E0B7    ;    //    lui x1 376366      ====        li ra, 0x5be2df00
                                                  30'd    5445    : data = 32'h    F0008093    ;    //    addi x1 x1 -256      ====        li ra, 0x5be2df00
                                                  30'd    5446    : data = 32'h    80000E37    ;    //    lui x28 524288      ====        li t3, 0x80000000
                                                  30'd    5447    : data = 32'h    000E0E13    ;    //    addi x28 x28 0      ====        li t3, 0x80000000
                                                  30'd    5448    : data = 32'h    DFECF097    ;    //    auipc x1 917199      ====        auipc ra, 917199
                                                  30'd    5449    : data = 32'h    ED179D97    ;    //    auipc x27 971129      ====        auipc s11, 971129
                                                  30'd    5450    : data = 32'h    DCD8BA97    ;    //    auipc x21 904587      ====        auipc s5, 904587
                                                  30'd    5451    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5452    : data = 32'h    65870A93    ;    //    addi x21 x14 1624      ====        addi s5, a4, 1624
                                                  30'd    5453    : data = 32'h    40E18A33    ;    //    sub x20 x3 x14      ====        sub s4, gp, a4
                                                  30'd    5454    : data = 32'h    395D8A13    ;    //    addi x20 x27 917      ====        addi s4, s11, 917
                                                  30'd    5455    : data = 32'h    011D8A33    ;    //    add x20 x27 x17      ====        add s4, s11, a7
                                                  30'd    5456    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5457    : data = 32'h    20170A13    ;    //    addi x20 x14 513      ====        addi s4, a4, 513
                                                  30'd    5458    : data = 32'h    F7AE4A97    ;    //    auipc x21 1014500      ====        auipc s5, 1014500
                                                  30'd    5459    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5460    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5461    : data = 32'h    34DE3A37    ;    //    lui x20 216547      ====        lui s4, 216547
                                                  30'd    5462    : data = 32'h    00840A33    ;    //    add x20 x8 x8      ====        add s4, s0, s0
                                                  30'd    5463    : data = 32'h    9185E417    ;    //    auipc x8 596062      ====        auipc s0, 596062
                                                  30'd    5464    : data = 32'h    EC6811B7    ;    //    lui x3 968321      ====        lui gp, 968321
                                                  30'd    5465    : data = 32'h    1D2E7437    ;    //    lui x8 119527      ====        lui s0, 119527
                                                  30'd    5466    : data = 32'h    331D8893    ;    //    addi x17 x27 817      ====        addi a7, s11, 817
                                                  30'd    5467    : data = 32'h    003881B3    ;    //    add x3 x17 x3      ====        add gp, a7, gp
                                                  30'd    5468    : data = 32'h    DB6A8093    ;    //    addi x1 x21 -586      ====        addi ra, s5, -586
                                                  30'd    5469    : data = 32'h    C54B9097    ;    //    auipc x1 808121      ====        auipc ra, 808121
                                                  30'd    5470    : data = 32'h    40210733    ;    //    sub x14 x2 x2      ====        sub a4, sp, sp
                                                  30'd    5471    : data = 32'h    01440133    ;    //    add x2 x8 x20      ====        add sp, s0, s4
                                                  30'd    5472    : data = 32'h    168060EF    ;    //    jal x1 24936      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_31
                                                  30'd    5473    : data = 32'h    01CA8FB3    ;    //    add x31 x21 x28      ====        add t6, s5, t3
                                                  30'd    5474    : data = 32'h    7ABC4913    ;    //    xori x18 x24 1963      ====        xori s2, s8, 1963
                                                  30'd    5475    : data = 32'h    86FA8D93    ;    //    addi x27 x21 -1937      ====        addi s11, s5, -1937
                                                  30'd    5476    : data = 32'h    54CBC593    ;    //    xori x11 x23 1356      ====        xori a1, s7, 1356
                                                  30'd    5477    : data = 32'h    016F9D33    ;    //    sll x26 x31 x22      ====        sll s10, t6, s6
                                                  30'd    5478    : data = 32'h    011958B3    ;    //    srl x17 x18 x17      ====        srl a7, s2, a7
                                                  30'd    5479    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5480    : data = 32'h    0087FCB3    ;    //    and x25 x15 x8      ====        and s9, a5, s0
                                                  30'd    5481    : data = 32'h    B564E993    ;    //    ori x19 x9 -1194      ====        ori s3, s1, -1194
                                                  30'd    5482    : data = 32'h    000CE033    ;    //    or x0 x25 x0      ====        or zero, s9, zero
                                                  30'd    5483    : data = 32'h    4165DCB3    ;    //    sra x25 x11 x22      ====        sra s9, a1, s6
                                                  30'd    5484    : data = 32'h    00AA9E93    ;    //    slli x29 x21 10      ====        slli t4, s5, 10
                                                  30'd    5485    : data = 32'h    0052E5B3    ;    //    or x11 x5 x5      ====        or a1, t0, t0
                                                  30'd    5486    : data = 32'h    0B243B13    ;    //    sltiu x22 x8 178      ====        sltiu s6, s0, 178
                                                  30'd    5487    : data = 32'h    010B8DB3    ;    //    add x27 x23 x16      ====        add s11, s7, a6
                                                  30'd    5488    : data = 32'h    D9678613    ;    //    addi x12 x15 -618      ====        addi a2, a5, -618
                                                  30'd    5489    : data = 32'h    01862D33    ;    //    slt x26 x12 x24      ====        slt s10, a2, s8
                                                  30'd    5490    : data = 32'h    01FAD7B3    ;    //    srl x15 x21 x31      ====        srl a5, s5, t6
                                                  30'd    5491    : data = 32'h    95AD1717    ;    //    auipc x14 613073      ====        auipc a4, 613073
                                                  30'd    5492    : data = 32'h    016E9A33    ;    //    sll x20 x29 x22      ====        sll s4, t4, s6
                                                  30'd    5493    : data = 32'h    01811813    ;    //    slli x16 x2 24      ====        slli a6, sp, 24
                                                  30'd    5494    : data = 32'h    000A7833    ;    //    and x16 x20 x0      ====        and a6, s4, zero
                                                  30'd    5495    : data = 32'h    40CF0B33    ;    //    sub x22 x30 x12      ====        sub s6, t5, a2
                                                  30'd    5496    : data = 32'h    309755B7    ;    //    lui x11 199029      ====        lui a1, 199029
                                                  30'd    5497    : data = 32'h    0088AB33    ;    //    slt x22 x17 x8      ====        slt s6, a7, s0
                                                  30'd    5498    : data = 32'h    7C96C813    ;    //    xori x16 x13 1993      ====        xori a6, a3, 1993
                                                  30'd    5499    : data = 32'h    F8E3A993    ;    //    slti x19 x7 -114      ====        slti s3, t2, -114
                                                  30'd    5500    : data = 32'h    007360B3    ;    //    or x1 x6 x7      ====        or ra, t1, t2
                                                  30'd    5501    : data = 32'h    01289E13    ;    //    slli x28 x17 18      ====        slli t3, a7, 18
                                                  30'd    5502    : data = 32'h    A1586893    ;    //    ori x17 x16 -1515      ====        ori a7, a6, -1515
                                                  30'd    5503    : data = 32'h    01045D13    ;    //    srli x26 x8 16      ====        srli s10, s0, 16
                                                  30'd    5504    : data = 32'h    77C57EB7    ;    //    lui x29 490583      ====        lui t4, 490583
                                                  30'd    5505    : data = 32'h    01461133    ;    //    sll x2 x12 x20      ====        sll sp, a2, s4
                                                  30'd    5506    : data = 32'h    014EC3B3    ;    //    xor x7 x29 x20      ====        xor t2, t4, s4
                                                  30'd    5507    : data = 32'h    5BF66093    ;    //    ori x1 x12 1471      ====        ori ra, a2, 1471
                                                  30'd    5508    : data = 32'h    01ABAC33    ;    //    slt x24 x23 x26      ====        slt s8, s7, s10
                                                  30'd    5509    : data = 32'h    01691AB3    ;    //    sll x21 x18 x22      ====        sll s5, s2, s6
                                                  30'd    5510    : data = 32'h    016D9333    ;    //    sll x6 x27 x22      ====        sll t1, s11, s6
                                                  30'd    5511    : data = 32'h    01F21C33    ;    //    sll x24 x4 x31      ====        sll s8, tp, t6
                                                  30'd    5512    : data = 32'h    01F85693    ;    //    srli x13 x16 31      ====        srli a3, a6, 31
                                                  30'd    5513    : data = 32'h    003341B3    ;    //    xor x3 x6 x3      ====        xor gp, t1, gp
                                                  30'd    5514    : data = 32'h    1A7D4813    ;    //    xori x16 x26 423      ====        xori a6, s10, 423
                                                  30'd    5515    : data = 32'h    2EFAA793    ;    //    slti x15 x21 751      ====        slti a5, s5, 751
                                                  30'd    5516    : data = 32'h    3D252613    ;    //    slti x12 x10 978      ====        slti a2, a0, 978
                                                  30'd    5517    : data = 32'h    72613637    ;    //    lui x12 468499      ====        lui a2, 468499
                                                  30'd    5518    : data = 32'h    029ACD13    ;    //    xori x26 x21 41      ====        xori s10, s5, 41
                                                  30'd    5519    : data = 32'h    018A9993    ;    //    slli x19 x21 24      ====        slli s3, s5, 24
                                                  30'd    5520    : data = 32'h    0188F833    ;    //    and x16 x17 x24      ====        and a6, a7, s8
                                                  30'd    5521    : data = 32'h    00824133    ;    //    xor x2 x4 x8      ====        xor sp, tp, s0
                                                  30'd    5522    : data = 32'h    00BBFDB3    ;    //    and x27 x23 x11      ====        and s11, s7, a1
                                                  30'd    5523    : data = 32'h    01724A33    ;    //    xor x20 x4 x23      ====        xor s4, tp, s7
                                                  30'd    5524    : data = 32'h    D54947B7    ;    //    lui x15 873620      ====        lui a5, 873620
                                                  30'd    5525    : data = 32'h    00762B33    ;    //    slt x22 x12 x7      ====        slt s6, a2, t2
                                                  30'd    5526    : data = 32'h    39DB6A13    ;    //    ori x20 x22 925      ====        ori s4, s6, 925
                                                  30'd    5527    : data = 32'h    41BB8FB3    ;    //    sub x31 x23 x27      ====        sub t6, s7, s11
                                                  30'd    5528    : data = 32'h    01D71CB3    ;    //    sll x25 x14 x29      ====        sll s9, a4, t4
                                                  30'd    5529    : data = 32'h    01D62FB3    ;    //    slt x31 x12 x29      ====        slt t6, a2, t4
                                                  30'd    5530    : data = 32'h    0135CA33    ;    //    xor x20 x11 x19      ====        xor s4, a1, s3
                                                  30'd    5531    : data = 32'h    FA4B4C37    ;    //    lui x24 1025204      ====        lui s8, 1025204
                                                  30'd    5532    : data = 32'h    01F409B3    ;    //    add x19 x8 x31      ====        add s3, s0, t6
                                                  30'd    5533    : data = 32'h    008C9AB3    ;    //    sll x21 x25 x8      ====        sll s5, s9, s0
                                                  30'd    5534    : data = 32'h    01BBF133    ;    //    and x2 x23 x27      ====        and sp, s7, s11
                                                  30'd    5535    : data = 32'h    000BA0B3    ;    //    slt x1 x23 x0      ====        slt ra, s7, zero
                                                  30'd    5536    : data = 32'h    01995E33    ;    //    srl x28 x18 x25      ====        srl t3, s2, s9
                                                  30'd    5537    : data = 32'h    001A6633    ;    //    or x12 x20 x1      ====        or a2, s4, ra
                                                  30'd    5538    : data = 32'h    B884CD13    ;    //    xori x26 x9 -1144      ====        xori s10, s1, -1144
                                                  30'd    5539    : data = 32'h    50B8AB93    ;    //    slti x23 x17 1291      ====        slti s7, a7, 1291
                                                  30'd    5540    : data = 32'h    00A7DFB3    ;    //    srl x31 x15 x10      ====        srl t6, a5, a0
                                                  30'd    5541    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5542    : data = 32'h    F5F10F93    ;    //    addi x31 x2 -161      ====        addi t6, sp, -161
                                                  30'd    5543    : data = 32'h    4186D313    ;    //    srai x6 x13 24      ====        srai t1, a3, 24
                                                  30'd    5544    : data = 32'h    40105E13    ;    //    srai x28 x0 1      ====        srai t3, zero, 1
                                                  30'd    5545    : data = 32'h    14AFB017    ;    //    auipc x0 84731      ====        auipc zero, 84731
                                                  30'd    5546    : data = 32'h    A0508293    ;    //    addi x5 x1 -1531      ====        addi t0, ra, -1531
                                                  30'd    5547    : data = 32'h    3A682E13    ;    //    slti x28 x16 934      ====        slti t3, a6, 934
                                                  30'd    5548    : data = 32'h    012DB8B3    ;    //    sltu x17 x27 x18      ====        sltu a7, s11, s2
                                                  30'd    5549    : data = 32'h    D6D5CD13    ;    //    xori x26 x11 -659      ====        xori s10, a1, -659
                                                  30'd    5550    : data = 32'h    3A3E4613    ;    //    xori x12 x28 931      ====        xori a2, t3, 931
                                                  30'd    5551    : data = 32'h    B1F34193    ;    //    xori x3 x6 -1249      ====        xori gp, t1, -1249
                                                  30'd    5552    : data = 32'h    00714833    ;    //    xor x16 x2 x7      ====        xor a6, sp, t2
                                                  30'd    5553    : data = 32'h    F28EEE93    ;    //    ori x29 x29 -216      ====        ori t4, t4, -216
                                                  30'd    5554    : data = 32'h    337DA137    ;    //    lui x2 210906      ====        lui sp, 210906
                                                  30'd    5555    : data = 32'h    01DC76B3    ;    //    and x13 x24 x29      ====        and a3, s8, t4
                                                  30'd    5556    : data = 32'h    005745B3    ;    //    xor x11 x14 x5      ====        xor a1, a4, t0
                                                  30'd    5557    : data = 32'h    71716E13    ;    //    ori x28 x2 1815      ====        ori t3, sp, 1815
                                                  30'd    5558    : data = 32'h    67670B93    ;    //    addi x23 x14 1654      ====        addi s7, a4, 1654
                                                  30'd    5559    : data = 32'h    41EC09B3    ;    //    sub x19 x24 x30      ====        sub s3, s8, t5
                                                  30'd    5560    : data = 32'h    56EA8A13    ;    //    addi x20 x21 1390      ====        addi s4, s5, 1390
                                                  30'd    5561    : data = 32'h    00F79E33    ;    //    sll x28 x15 x15      ====        sll t3, a5, a5
                                                  30'd    5562    : data = 32'h    010338B3    ;    //    sltu x17 x6 x16      ====        sltu a7, t1, a6
                                                  30'd    5563    : data = 32'h    01B867B3    ;    //    or x15 x16 x27      ====        or a5, a6, s11
                                                  30'd    5564    : data = 32'h    8E354A93    ;    //    xori x21 x10 -1821      ====        xori s5, a0, -1821
                                                  30'd    5565    : data = 32'h    68043593    ;    //    sltiu x11 x8 1664      ====        sltiu a1, s0, 1664
                                                  30'd    5566    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5567    : data = 32'h    01C93733    ;    //    sltu x14 x18 x28      ====        sltu a4, s2, t3
                                                  30'd    5568    : data = 32'h    40800733    ;    //    sub x14 x0 x8      ====        sub a4, zero, s0
                                                  30'd    5569    : data = 32'h    D96157B7    ;    //    lui x15 890389      ====        lui a5, 890389
                                                  30'd    5570    : data = 32'h    01A21433    ;    //    sll x8 x4 x26      ====        sll s0, tp, s10
                                                  30'd    5571    : data = 32'h    01CE1D33    ;    //    sll x26 x28 x28      ====        sll s10, t3, t3
                                                  30'd    5572    : data = 32'h    00BDD893    ;    //    srli x17 x27 11      ====        srli a7, s11, 11
                                                  30'd    5573    : data = 32'h    0082E733    ;    //    or x14 x5 x8      ====        or a4, t0, s0
                                                  30'd    5574    : data = 32'h    00DC5BB3    ;    //    srl x23 x24 x13      ====        srl s7, s8, a3
                                                  30'd    5575    : data = 32'h    6665B493    ;    //    sltiu x9 x11 1638      ====        sltiu s1, a1, 1638
                                                  30'd    5576    : data = 32'h    16132D13    ;    //    slti x26 x6 353      ====        slti s10, t1, 353
                                                  30'd    5577    : data = 32'h    40688333    ;    //    sub x6 x17 x6      ====        sub t1, a7, t1
                                                  30'd    5578    : data = 32'h    00C9F033    ;    //    and x0 x19 x12      ====        and zero, s3, a2
                                                  30'd    5579    : data = 32'h    01D2DC93    ;    //    srli x25 x5 29      ====        srli s9, t0, 29
                                                  30'd    5580    : data = 32'h    2F6F3D17    ;    //    auipc x26 194291      ====        auipc s10, 194291
                                                  30'd    5581    : data = 32'h    014D1793    ;    //    slli x15 x26 20      ====        slli a5, s10, 20
                                                  30'd    5582    : data = 32'h    01C51993    ;    //    slli x19 x10 28      ====        slli s3, a0, 28
                                                  30'd    5583    : data = 32'h    17EFFD13    ;    //    andi x26 x31 382      ====        andi s10, t6, 382
                                                  30'd    5584    : data = 32'h    405F5FB3    ;    //    sra x31 x30 x5      ====        sra t6, t5, t0
                                                  30'd    5585    : data = 32'h    012FA2B3    ;    //    slt x5 x31 x18      ====        slt t0, t6, s2
                                                  30'd    5586    : data = 32'h    A5A73137    ;    //    lui x2 678515      ====        lui sp, 678515
                                                  30'd    5587    : data = 32'h    0144DBB3    ;    //    srl x23 x9 x20      ====        srl s7, s1, s4
                                                  30'd    5588    : data = 32'h    41FF52B3    ;    //    sra x5 x30 x31      ====        sra t0, t5, t6
                                                  30'd    5589    : data = 32'h    5D53B913    ;    //    sltiu x18 x7 1493      ====        sltiu s2, t2, 1493
                                                  30'd    5590    : data = 32'h    012340B3    ;    //    xor x1 x6 x18      ====        xor ra, t1, s2
                                                  30'd    5591    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5592    : data = 32'h    014F74B3    ;    //    and x9 x30 x20      ====        and s1, t5, s4
                                                  30'd    5593    : data = 32'h    01C91413    ;    //    slli x8 x18 28      ====        slli s0, s2, 28
                                                  30'd    5594    : data = 32'h    0070FEB3    ;    //    and x29 x1 x7      ====        and t4, ra, t2
                                                  30'd    5595    : data = 32'h    DD4E6D13    ;    //    ori x26 x28 -556      ====        ori s10, t3, -556
                                                  30'd    5596    : data = 32'h    2E4F6E13    ;    //    ori x28 x30 740      ====        ori t3, t5, 740
                                                  30'd    5597    : data = 32'h    409255B3    ;    //    sra x11 x4 x9      ====        sra a1, tp, s1
                                                  30'd    5598    : data = 32'h    008207B3    ;    //    add x15 x4 x8      ====        add a5, tp, s0
                                                  30'd    5599    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5600    : data = 32'h    3E99DE37    ;    //    lui x28 256413      ====        lui t3, 256413
                                                  30'd    5601    : data = 32'h    99EFC993    ;    //    xori x19 x31 -1634      ====        xori s3, t6, -1634
                                                  30'd    5602    : data = 32'h    41CC54B3    ;    //    sra x9 x24 x28      ====        sra s1, s8, t3
                                                  30'd    5603    : data = 32'h    4162DE93    ;    //    srai x29 x5 22      ====        srai t4, t0, 22
                                                  30'd    5604    : data = 32'h    01F7DA13    ;    //    srli x20 x15 31      ====        srli s4, a5, 31
                                                  30'd    5605    : data = 32'h    00049CB3    ;    //    sll x25 x9 x0      ====        sll s9, s1, zero
                                                  30'd    5606    : data = 32'h    00C0A6B3    ;    //    slt x13 x1 x12      ====        slt a3, ra, a2
                                                  30'd    5607    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5608    : data = 32'h    00BD0733    ;    //    add x14 x26 x11      ====        add a4, s10, a1
                                                  30'd    5609    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5610    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5611    : data = 32'h    015011B3    ;    //    sll x3 x0 x21      ====        sll gp, zero, s5
                                                  30'd    5612    : data = 32'h    F3001B37    ;    //    lui x22 995329      ====        lui s6, 995329
                                                  30'd    5613    : data = 32'h    D9627A13    ;    //    andi x20 x4 -618      ====        andi s4, tp, -618
                                                  30'd    5614    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5615    : data = 32'h    402ED713    ;    //    srai x14 x29 2      ====        srai a4, t4, 2
                                                  30'd    5616    : data = 32'h    01DFD813    ;    //    srli x16 x31 29      ====        srli a6, t6, 29
                                                  30'd    5617    : data = 32'h    3018C413    ;    //    xori x8 x17 769      ====        xori s0, a7, 769
                                                  30'd    5618    : data = 32'h    00671CB3    ;    //    sll x25 x14 x6      ====        sll s9, a4, t1
                                                  30'd    5619    : data = 32'h    E2623613    ;    //    sltiu x12 x4 -474      ====        sltiu a2, tp, -474
                                                  30'd    5620    : data = 32'h    00BBC933    ;    //    xor x18 x23 x11      ====        xor s2, s7, a1
                                                  30'd    5621    : data = 32'h    0EDE0597    ;    //    auipc x11 60896      ====        auipc a1, 60896
                                                  30'd    5622    : data = 32'h    013C1693    ;    //    slli x13 x24 19      ====        slli a3, s8, 19
                                                  30'd    5623    : data = 32'h    004D92B3    ;    //    sll x5 x27 x4      ====        sll t0, s11, tp
                                                  30'd    5624    : data = 32'h    41CFDEB3    ;    //    sra x29 x31 x28      ====        sra t4, t6, t3
                                                  30'd    5625    : data = 32'h    24E15317    ;    //    auipc x6 151061      ====        auipc t1, 151061
                                                  30'd    5626    : data = 32'h    01E7EA33    ;    //    or x20 x15 x30      ====        or s4, a5, t5
                                                  30'd    5627    : data = 32'h    7095A4B7    ;    //    lui x9 461146      ====        lui s1, 461146
                                                  30'd    5628    : data = 32'h    DD8467B7    ;    //    lui x15 907334      ====        lui a5, 907334
                                                  30'd    5629    : data = 32'h    00DCE4B3    ;    //    or x9 x25 x13      ====        or s1, s9, a3
                                                  30'd    5630    : data = 32'h    1674E693    ;    //    ori x13 x9 359      ====        ori a3, s1, 359
                                                  30'd    5631    : data = 32'h    D31D7317    ;    //    auipc x6 864727      ====        auipc t1, 864727
                                                  30'd    5632    : data = 32'h    170E8613    ;    //    addi x12 x29 368      ====        addi a2, t4, 368
                                                  30'd    5633    : data = 32'h    415153B3    ;    //    sra x7 x2 x21      ====        sra t2, sp, s5
                                                  30'd    5634    : data = 32'h    38AB5637    ;    //    lui x12 232117      ====        lui a2, 232117
                                                  30'd    5635    : data = 32'h    62D2CF93    ;    //    xori x31 x5 1581      ====        xori t6, t0, 1581
                                                  30'd    5636    : data = 32'h    005FCD33    ;    //    xor x26 x31 x5      ====        xor s10, t6, t0
                                                  30'd    5637    : data = 32'h    FEA4B817    ;    //    auipc x16 1043019      ====        auipc a6, 1043019
                                                  30'd    5638    : data = 32'h    2FAF2813    ;    //    slti x16 x30 762      ====        slti a6, t5, 762
                                                  30'd    5639    : data = 32'h    019DEBB3    ;    //    or x23 x27 x25      ====        or s7, s11, s9
                                                  30'd    5640    : data = 32'h    00AF1733    ;    //    sll x14 x30 x10      ====        sll a4, t5, a0
                                                  30'd    5641    : data = 32'h    412DD313    ;    //    srai x6 x27 18      ====        srai t1, s11, 18
                                                  30'd    5642    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5643    : data = 32'h    01D0C833    ;    //    xor x16 x1 x29      ====        xor a6, ra, t4
                                                  30'd    5644    : data = 32'h    37696613    ;    //    ori x12 x18 886      ====        ori a2, s2, 886
                                                  30'd    5645    : data = 32'h    004F9913    ;    //    slli x18 x31 4      ====        slli s2, t6, 4
                                                  30'd    5646    : data = 32'h    00F45DB3    ;    //    srl x27 x8 x15      ====        srl s11, s0, a5
                                                  30'd    5647    : data = 32'h    01FBAEB3    ;    //    slt x29 x23 x31      ====        slt t4, s7, t6
                                                  30'd    5648    : data = 32'h    9828ED93    ;    //    ori x27 x17 -1662      ====        ori s11, a7, -1662
                                                  30'd    5649    : data = 32'h    FD6A0993    ;    //    addi x19 x20 -42      ====        addi s3, s4, -42
                                                  30'd    5650    : data = 32'h    00ED5A93    ;    //    srli x21 x26 14      ====        srli s5, s10, 14
                                                  30'd    5651    : data = 32'h    40045FB3    ;    //    sra x31 x8 x0      ====        sra t6, s0, zero
                                                  30'd    5652    : data = 32'h    2760F413    ;    //    andi x8 x1 630      ====        andi s0, ra, 630
                                                  30'd    5653    : data = 32'h    00EA7633    ;    //    and x12 x20 x14      ====        and a2, s4, a4
                                                  30'd    5654    : data = 32'h    00F5ADB3    ;    //    slt x27 x11 x15      ====        slt s11, a1, a5
                                                  30'd    5655    : data = 32'h    92092E13    ;    //    slti x28 x18 -1760      ====        slti t3, s2, -1760
                                                  30'd    5656    : data = 32'h    4D203413    ;    //    sltiu x8 x0 1234      ====        sltiu s0, zero, 1234
                                                  30'd    5657    : data = 32'h    01F61433    ;    //    sll x8 x12 x31      ====        sll s0, a2, t6
                                                  30'd    5658    : data = 32'h    019F40B3    ;    //    xor x1 x30 x25      ====        xor ra, t5, s9
                                                  30'd    5659    : data = 32'h    4151DB93    ;    //    srai x23 x3 21      ====        srai s7, gp, 21
                                                  30'd    5660    : data = 32'h    CC262B93    ;    //    slti x23 x12 -830      ====        slti s7, a2, -830
                                                  30'd    5661    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5662    : data = 32'h    00D8CBB3    ;    //    xor x23 x17 x13      ====        xor s7, a7, a3
                                                  30'd    5663    : data = 32'h    019CD333    ;    //    srl x6 x25 x25      ====        srl t1, s9, s9
                                                  30'd    5664    : data = 32'h    014090B3    ;    //    sll x1 x1 x20      ====        sll ra, ra, s4
                                                  30'd    5665    : data = 32'h    001EECB3    ;    //    or x25 x29 x1      ====        or s9, t4, ra
                                                  30'd    5666    : data = 32'h    7CA6E013    ;    //    ori x0 x13 1994      ====        ori zero, a3, 1994
                                                  30'd    5667    : data = 32'h    019FB333    ;    //    sltu x6 x31 x25      ====        sltu t1, t6, s9
                                                  30'd    5668    : data = 32'h    01C0D033    ;    //    srl x0 x1 x28      ====        srl zero, ra, t3
                                                  30'd    5669    : data = 32'h    015AFA33    ;    //    and x20 x21 x21      ====        and s4, s5, s5
                                                  30'd    5670    : data = 32'h    00AED9B3    ;    //    srl x19 x29 x10      ====        srl s3, t4, a0
                                                  30'd    5671    : data = 32'h    0008DA93    ;    //    srli x21 x17 0      ====        srli s5, a7, 0
                                                  30'd    5672    : data = 32'h    83714497    ;    //    auipc x9 538388      ====        auipc s1, 538388
                                                  30'd    5673    : data = 32'h    01439E33    ;    //    sll x28 x7 x20      ====        sll t3, t2, s4
                                                  30'd    5674    : data = 32'h    00229313    ;    //    slli x6 x5 2      ====        slli t1, t0, 2
                                                  30'd    5675    : data = 32'h    B2D695B7    ;    //    lui x11 732521      ====        lui a1, 732521
                                                  30'd    5676    : data = 32'h    50D49897    ;    //    auipc x17 331081      ====        auipc a7, 331081
                                                  30'd    5677    : data = 32'h    B3E878B7    ;    //    lui x17 736903      ====        lui a7, 736903
                                                  30'd    5678    : data = 32'h    07284893    ;    //    xori x17 x16 114      ====        xori a7, a6, 114
                                                  30'd    5679    : data = 32'h    9C8841B7    ;    //    lui x3 641156      ====        lui gp, 641156
                                                  30'd    5680    : data = 32'h    01AC62B3    ;    //    or x5 x24 x26      ====        or t0, s8, s10
                                                  30'd    5681    : data = 32'h    3390A693    ;    //    slti x13 x1 825      ====        slti a3, ra, 825
                                                  30'd    5682    : data = 32'h    0038F2B3    ;    //    and x5 x17 x3      ====        and t0, a7, gp
                                                  30'd    5683    : data = 32'h    000DD013    ;    //    srli x0 x27 0      ====        srli zero, s11, 0
                                                  30'd    5684    : data = 32'h    EB1EC013    ;    //    xori x0 x29 -335      ====        xori zero, t4, -335
                                                  30'd    5685    : data = 32'h    4160D913    ;    //    srai x18 x1 22      ====        srai s2, ra, 22
                                                  30'd    5686    : data = 32'h    4C5A3313    ;    //    sltiu x6 x20 1221      ====        sltiu t1, s4, 1221
                                                  30'd    5687    : data = 32'h    405A82B3    ;    //    sub x5 x21 x5      ====        sub t0, s5, t0
                                                  30'd    5688    : data = 32'h    015B7133    ;    //    and x2 x22 x21      ====        and sp, s6, s5
                                                  30'd    5689    : data = 32'h    00CB6A33    ;    //    or x20 x22 x12      ====        or s4, s6, a2
                                                  30'd    5690    : data = 32'h    01EF6833    ;    //    or x16 x30 x30      ====        or a6, t5, t5
                                                  30'd    5691    : data = 32'h    89BB6FB7    ;    //    lui x31 564150      ====        lui t6, 564150
                                                  30'd    5692    : data = 32'h    B6C67013    ;    //    andi x0 x12 -1172      ====        andi zero, a2, -1172
                                                  30'd    5693    : data = 32'h    00E055B3    ;    //    srl x11 x0 x14      ====        srl a1, zero, a4
                                                  30'd    5694    : data = 32'h    0010EAB3    ;    //    or x21 x1 x1      ====        or s5, ra, ra
                                                  30'd    5695    : data = 32'h    01CD5413    ;    //    srli x8 x26 28      ====        srli s0, s10, 28
                                                  30'd    5696    : data = 32'h    78C86693    ;    //    ori x13 x16 1932      ====        ori a3, a6, 1932
                                                  30'd    5697    : data = 32'h    A9594637    ;    //    lui x12 693652      ====        lui a2, 693652
                                                  30'd    5698    : data = 32'h    01E69593    ;    //    slli x11 x13 30      ====        slli a1, a3, 30
                                                  30'd    5699    : data = 32'h    00611813    ;    //    slli x16 x2 6      ====        slli a6, sp, 6
                                                  30'd    5700    : data = 32'h    00D86EB3    ;    //    or x29 x16 x13      ====        or t4, a6, a3
                                                  30'd    5701    : data = 32'h    4058D893    ;    //    srai x17 x17 5      ====        srai a7, a7, 5
                                                  30'd    5702    : data = 32'h    9234F4B7    ;    //    lui x9 598863      ====        lui s1, 598863
                                                  30'd    5703    : data = 32'h    41A28DB3    ;    //    sub x27 x5 x26      ====        sub s11, t0, s10
                                                  30'd    5704    : data = 32'h    00FC0133    ;    //    add x2 x24 x15      ====        add sp, s8, a5
                                                  30'd    5705    : data = 32'h    01A7AAB3    ;    //    slt x21 x15 x26      ====        slt s5, a5, s10
                                                  30'd    5706    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5707    : data = 32'h    F4896917    ;    //    auipc x18 1001622      ====        auipc s2, 1001622
                                                  30'd    5708    : data = 32'h    58FD2713    ;    //    slti x14 x26 1423      ====        slti a4, s10, 1423
                                                  30'd    5709    : data = 32'h    41215893    ;    //    srai x17 x2 18      ====        srai a7, sp, 18
                                                  30'd    5710    : data = 32'h    0194E833    ;    //    or x16 x9 x25      ====        or a6, s1, s9
                                                  30'd    5711    : data = 32'h    41878333    ;    //    sub x6 x15 x24      ====        sub t1, a5, s8
                                                  30'd    5712    : data = 32'h    00501D93    ;    //    slli x27 x0 5      ====        slli s11, zero, 5
                                                  30'd    5713    : data = 32'h    00468B33    ;    //    add x22 x13 x4      ====        add s6, a3, tp
                                                  30'd    5714    : data = 32'h    00B6BE33    ;    //    sltu x28 x13 x11      ====        sltu t3, a3, a1
                                                  30'd    5715    : data = 32'h    84A1E613    ;    //    ori x12 x3 -1974      ====        ori a2, gp, -1974
                                                  30'd    5716    : data = 32'h    A996A193    ;    //    slti x3 x13 -1383      ====        slti gp, a3, -1383
                                                  30'd    5717    : data = 32'h    40F85F93    ;    //    srai x31 x16 15      ====        srai t6, a6, 15
                                                  30'd    5718    : data = 32'h    401384B3    ;    //    sub x9 x7 x1      ====        sub s1, t2, ra
                                                  30'd    5719    : data = 32'h    E017AD93    ;    //    slti x27 x15 -511      ====        slti s11, a5, -511
                                                  30'd    5720    : data = 32'h    27C05BB7    ;    //    lui x23 162821      ====        lui s7, 162821
                                                  30'd    5721    : data = 32'h    01B3E833    ;    //    or x16 x7 x27      ====        or a6, t2, s11
                                                  30'd    5722    : data = 32'h    405650B3    ;    //    sra x1 x12 x5      ====        sra ra, a2, t0
                                                  30'd    5723    : data = 32'h    01C51F93    ;    //    slli x31 x10 28      ====        slli t6, a0, 28
                                                  30'd    5724    : data = 32'h    5552F493    ;    //    andi x9 x5 1365      ====        andi s1, t0, 1365
                                                  30'd    5725    : data = 32'h    01BAAE33    ;    //    slt x28 x21 x27      ====        slt t3, s5, s11
                                                  30'd    5726    : data = 32'h    208BBDB7    ;    //    lui x27 133307      ====        lui s11, 133307
                                                  30'd    5727    : data = 32'h    017B1833    ;    //    sll x16 x22 x23      ====        sll a6, s6, s7
                                                  30'd    5728    : data = 32'h    89F58813    ;    //    addi x16 x11 -1889      ====        addi a6, a1, -1889
                                                  30'd    5729    : data = 32'h    16C6B813    ;    //    sltiu x16 x13 364      ====        sltiu a6, a3, 364
                                                  30'd    5730    : data = 32'h    1A909317    ;    //    auipc x6 108809      ====        auipc t1, 108809
                                                  30'd    5731    : data = 32'h    01293633    ;    //    sltu x12 x18 x18      ====        sltu a2, s2, s2
                                                  30'd    5732    : data = 32'h    292B1717    ;    //    auipc x14 168625      ====        auipc a4, 168625
                                                  30'd    5733    : data = 32'h    00E2AFB3    ;    //    slt x31 x5 x14      ====        slt t6, t0, a4
                                                  30'd    5734    : data = 32'h    6C325717    ;    //    auipc x14 443173      ====        auipc a4, 443173
                                                  30'd    5735    : data = 32'h    DC4F2B93    ;    //    slti x23 x30 -572      ====        slti s7, t5, -572
                                                  30'd    5736    : data = 32'h    01EB9D13    ;    //    slli x26 x23 30      ====        slli s10, s7, 30
                                                  30'd    5737    : data = 32'h    783DB493    ;    //    sltiu x9 x27 1923      ====        sltiu s1, s11, 1923
                                                  30'd    5738    : data = 32'h    010742B3    ;    //    xor x5 x14 x16      ====        xor t0, a4, a6
                                                  30'd    5739    : data = 32'h    0026D5B3    ;    //    srl x11 x13 x2      ====        srl a1, a3, sp
                                                  30'd    5740    : data = 32'h    0129B1B3    ;    //    sltu x3 x19 x18      ====        sltu gp, s3, s2
                                                  30'd    5741    : data = 32'h    009BC033    ;    //    xor x0 x23 x9      ====        xor zero, s7, s1
                                                  30'd    5742    : data = 32'h    411D51B3    ;    //    sra x3 x26 x17      ====        sra gp, s10, a7
                                                  30'd    5743    : data = 32'h    018A1593    ;    //    slli x11 x20 24      ====        slli a1, s4, 24
                                                  30'd    5744    : data = 32'h    8D277613    ;    //    andi x12 x14 -1838      ====        andi a2, a4, -1838
                                                  30'd    5745    : data = 32'h    406F52B3    ;    //    sra x5 x30 x6      ====        sra t0, t5, t1
                                                  30'd    5746    : data = 32'h    8C8F3D93    ;    //    sltiu x27 x30 -1848      ====        sltiu s11, t5, -1848
                                                  30'd    5747    : data = 32'h    A9554693    ;    //    xori x13 x10 -1387      ====        xori a3, a0, -1387
                                                  30'd    5748    : data = 32'h    3E50E713    ;    //    ori x14 x1 997      ====        ori a4, ra, 997
                                                  30'd    5749    : data = 32'h    77637F93    ;    //    andi x31 x6 1910      ====        andi t6, t1, 1910
                                                  30'd    5750    : data = 32'h    40175F93    ;    //    srai x31 x14 1      ====        srai t6, a4, 1
                                                  30'd    5751    : data = 32'h    4100D6B3    ;    //    sra x13 x1 x16      ====        sra a3, ra, a6
                                                  30'd    5752    : data = 32'h    00BF64B3    ;    //    or x9 x30 x11      ====        or s1, t5, a1
                                                  30'd    5753    : data = 32'h    00191D33    ;    //    sll x26 x18 x1      ====        sll s10, s2, ra
                                                  30'd    5754    : data = 32'h    00B04AB3    ;    //    xor x21 x0 x11      ====        xor s5, zero, a1
                                                  30'd    5755    : data = 32'h    90ED1737    ;    //    lui x14 593617      ====        lui a4, 593617
                                                  30'd    5756    : data = 32'h    008AD713    ;    //    srli x14 x21 8      ====        srli a4, s5, 8
                                                  30'd    5757    : data = 32'h    40160433    ;    //    sub x8 x12 x1      ====        sub s0, a2, ra
                                                  30'd    5758    : data = 32'h    B7F50B13    ;    //    addi x22 x10 -1153      ====        addi s6, a0, -1153
                                                  30'd    5759    : data = 32'h    01507933    ;    //    and x18 x0 x21      ====        and s2, zero, s5
                                                  30'd    5760    : data = 32'h    4FFF7C13    ;    //    andi x24 x30 1279      ====        andi s8, t5, 1279
                                                  30'd    5761    : data = 32'h    1E2A0093    ;    //    addi x1 x20 482      ====        addi ra, s4, 482
                                                  30'd    5762    : data = 32'h    0165B033    ;    //    sltu x0 x11 x22      ====        sltu zero, a1, s6
                                                  30'd    5763    : data = 32'h    AB1B0D13    ;    //    addi x26 x22 -1359      ====        addi s10, s6, -1359
                                                  30'd    5764    : data = 32'h    62D83013    ;    //    sltiu x0 x16 1581      ====        sltiu zero, a6, 1581
                                                  30'd    5765    : data = 32'h    003A3733    ;    //    sltu x14 x20 x3      ====        sltu a4, s4, gp
                                                  30'd    5766    : data = 32'h    4A66C113    ;    //    xori x2 x13 1190      ====        xori sp, a3, 1190
                                                  30'd    5767    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5768    : data = 32'h    013F72B3    ;    //    and x5 x30 x19      ====        and t0, t5, s3
                                                  30'd    5769    : data = 32'h    010B34B3    ;    //    sltu x9 x22 x16      ====        sltu s1, s6, a6
                                                  30'd    5770    : data = 32'h    41848633    ;    //    sub x12 x9 x24      ====        sub a2, s1, s8
                                                  30'd    5771    : data = 32'h    003515B3    ;    //    sll x11 x10 x3      ====        sll a1, a0, gp
                                                  30'd    5772    : data = 32'h    FF51BD13    ;    //    sltiu x26 x3 -11      ====        sltiu s10, gp, -11
                                                  30'd    5773    : data = 32'h    01EFFFB3    ;    //    and x31 x31 x30      ====        and t6, t6, t5
                                                  30'd    5774    : data = 32'h    007790B3    ;    //    sll x1 x15 x7      ====        sll ra, a5, t2
                                                  30'd    5775    : data = 32'h    B3EE4593    ;    //    xori x11 x28 -1218      ====        xori a1, t3, -1218
                                                  30'd    5776    : data = 32'h    30A80313    ;    //    addi x6 x16 778      ====        addi t1, a6, 778
                                                  30'd    5777    : data = 32'h    F49DC837    ;    //    lui x16 1001948      ====        lui a6, 1001948
                                                  30'd    5778    : data = 32'h    95CDCE13    ;    //    xori x28 x27 -1700      ====        xori t3, s11, -1700
                                                  30'd    5779    : data = 32'h    00623EB3    ;    //    sltu x29 x4 x6      ====        sltu t4, tp, t1
                                                  30'd    5780    : data = 32'h    008AA5B3    ;    //    slt x11 x21 x8      ====        slt a1, s5, s0
                                                  30'd    5781    : data = 32'h    E788AF93    ;    //    slti x31 x17 -392      ====        slti t6, a7, -392
                                                  30'd    5782    : data = 32'h    A3378E97    ;    //    auipc x29 668536      ====        auipc t4, 668536
                                                  30'd    5783    : data = 32'h    00CE4933    ;    //    xor x18 x28 x12      ====        xor s2, t3, a2
                                                  30'd    5784    : data = 32'h    AFE27E93    ;    //    andi x29 x4 -1282      ====        andi t4, tp, -1282
                                                  30'd    5785    : data = 32'h    019597B3    ;    //    sll x15 x11 x25      ====        sll a5, a1, s9
                                                  30'd    5786    : data = 32'h    006CA9B3    ;    //    slt x19 x25 x6      ====        slt s3, s9, t1
                                                  30'd    5787    : data = 32'h    011B5C33    ;    //    srl x24 x22 x17      ====        srl s8, s6, a7
                                                  30'd    5788    : data = 32'h    013884B3    ;    //    add x9 x17 x19      ====        add s1, a7, s3
                                                  30'd    5789    : data = 32'h    006B1A33    ;    //    sll x20 x22 x6      ====        sll s4, s6, t1
                                                  30'd    5790    : data = 32'h    80D14D13    ;    //    xori x26 x2 -2035      ====        xori s10, sp, -2035
                                                  30'd    5791    : data = 32'h    41FF8133    ;    //    sub x2 x31 x31      ====        sub sp, t6, t6
                                                  30'd    5792    : data = 32'h    8DB4C0B7    ;    //    lui x1 580428      ====        lui ra, 580428
                                                  30'd    5793    : data = 32'h    3B6F8893    ;    //    addi x17 x31 950      ====        addi a7, t6, 950
                                                  30'd    5794    : data = 32'h    019B1293    ;    //    slli x5 x22 25      ====        slli t0, s6, 25
                                                  30'd    5795    : data = 32'h    2D498713    ;    //    addi x14 x19 724      ====        addi a4, s3, 724
                                                  30'd    5796    : data = 32'h    011BD893    ;    //    srli x17 x23 17      ====        srli a7, s7, 17
                                                  30'd    5797    : data = 32'h    002C2A33    ;    //    slt x20 x24 x2      ====        slt s4, s8, sp
                                                  30'd    5798    : data = 32'h    01B697B3    ;    //    sll x15 x13 x27      ====        sll a5, a3, s11
                                                  30'd    5799    : data = 32'h    BE637713    ;    //    andi x14 x6 -1050      ====        andi a4, t1, -1050
                                                  30'd    5800    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5801    : data = 32'h    405350B3    ;    //    sra x1 x6 x5      ====        sra ra, t1, t0
                                                  30'd    5802    : data = 32'h    000A1A93    ;    //    slli x21 x20 0      ====        slli s5, s4, 0
                                                  30'd    5803    : data = 32'h    405B0133    ;    //    sub x2 x22 x5      ====        sub sp, s6, t0
                                                  30'd    5804    : data = 32'h    0080D413    ;    //    srli x8 x1 8      ====        srli s0, ra, 8
                                                  30'd    5805    : data = 32'h    00A84733    ;    //    xor x14 x16 x10      ====        xor a4, a6, a0
                                                  30'd    5806    : data = 32'h    0105A1B3    ;    //    slt x3 x11 x16      ====        slt gp, a1, a6
                                                  30'd    5807    : data = 32'h    0075BCB3    ;    //    sltu x25 x11 x7      ====        sltu s9, a1, t2
                                                  30'd    5808    : data = 32'h    31C86613    ;    //    ori x12 x16 796      ====        ori a2, a6, 796
                                                  30'd    5809    : data = 32'h    5AD7A1B7    ;    //    lui x3 372090      ====        lui gp, 372090
                                                  30'd    5810    : data = 32'h    E5302B13    ;    //    slti x22 x0 -429      ====        slti s6, zero, -429
                                                  30'd    5811    : data = 32'h    F4030093    ;    //    addi x1 x6 -192      ====        addi ra, t1, -192
                                                  30'd    5812    : data = 32'h    002D4AB3    ;    //    xor x21 x26 x2      ====        xor s5, s10, sp
                                                  30'd    5813    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5814    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5815    : data = 32'h    0109A433    ;    //    slt x8 x19 x16      ====        slt s0, s3, a6
                                                  30'd    5816    : data = 32'h    D66DCA13    ;    //    xori x20 x27 -666      ====        xori s4, s11, -666
                                                  30'd    5817    : data = 32'h    41A75FB3    ;    //    sra x31 x14 x26      ====        sra t6, a4, s10
                                                  30'd    5818    : data = 32'h    016436B3    ;    //    sltu x13 x8 x22      ====        sltu a3, s0, s6
                                                  30'd    5819    : data = 32'h    22A7F993    ;    //    andi x19 x15 554      ====        andi s3, a5, 554
                                                  30'd    5820    : data = 32'h    00E0C833    ;    //    xor x16 x1 x14      ====        xor a6, ra, a4
                                                  30'd    5821    : data = 32'h    00EA6633    ;    //    or x12 x20 x14      ====        or a2, s4, a4
                                                  30'd    5822    : data = 32'h    004F72B3    ;    //    and x5 x30 x4      ====        and t0, t5, tp
                                                  30'd    5823    : data = 32'h    3E022613    ;    //    slti x12 x4 992      ====        slti a2, tp, 992
                                                  30'd    5824    : data = 32'h    0171CD33    ;    //    xor x26 x3 x23      ====        xor s10, gp, s7
                                                  30'd    5825    : data = 32'h    3709A2B7    ;    //    lui x5 225434      ====        lui t0, 225434
                                                  30'd    5826    : data = 32'h    41110733    ;    //    sub x14 x2 x17      ====        sub a4, sp, a7
                                                  30'd    5827    : data = 32'h    41A70C93    ;    //    addi x25 x14 1050      ====        addi s9, a4, 1050
                                                  30'd    5828    : data = 32'h    40480AB3    ;    //    sub x21 x16 x4      ====        sub s5, a6, tp
                                                  30'd    5829    : data = 32'h    D4776113    ;    //    ori x2 x14 -697      ====        ori sp, a4, -697
                                                  30'd    5830    : data = 32'h    BB821C97    ;    //    auipc x25 768033      ====        auipc s9, 768033
                                                  30'd    5831    : data = 32'h    01269013    ;    //    slli x0 x13 18      ====        slli zero, a3, 18
                                                  30'd    5832    : data = 32'h    41F1DA13    ;    //    srai x20 x3 31      ====        srai s4, gp, 31
                                                  30'd    5833    : data = 32'h    41BB5C93    ;    //    srai x25 x22 27      ====        srai s9, s6, 27
                                                  30'd    5834    : data = 32'h    00714433    ;    //    xor x8 x2 x7      ====        xor s0, sp, t2
                                                  30'd    5835    : data = 32'h    0103DCB3    ;    //    srl x25 x7 x16      ====        srl s9, t2, a6
                                                  30'd    5836    : data = 32'h    A94C0397    ;    //    auipc x7 693440      ====        auipc t2, 693440
                                                  30'd    5837    : data = 32'h    B78A48B7    ;    //    lui x17 751780      ====        lui a7, 751780
                                                  30'd    5838    : data = 32'h    53C3E813    ;    //    ori x16 x7 1340      ====        ori a6, t2, 1340
                                                  30'd    5839    : data = 32'h    41B4D1B3    ;    //    sra x3 x9 x27      ====        sra gp, s1, s11
                                                  30'd    5840    : data = 32'h    AE330D37    ;    //    lui x26 713520      ====        lui s10, 713520
                                                  30'd    5841    : data = 32'h    9BC72D13    ;    //    slti x26 x14 -1604      ====        slti s10, a4, -1604
                                                  30'd    5842    : data = 32'h    00C3D8B3    ;    //    srl x17 x7 x12      ====        srl a7, t2, a2
                                                  30'd    5843    : data = 32'h    08D8F613    ;    //    andi x12 x17 141      ====        andi a2, a7, 141
                                                  30'd    5844    : data = 32'h    00864333    ;    //    xor x6 x12 x8      ====        xor t1, a2, s0
                                                  30'd    5845    : data = 32'h    E3DBA193    ;    //    slti x3 x23 -451      ====        slti gp, s7, -451
                                                  30'd    5846    : data = 32'h    40DA5313    ;    //    srai x6 x20 13      ====        srai t1, s4, 13
                                                  30'd    5847    : data = 32'h    F34AA337    ;    //    lui x6 996522      ====        lui t1, 996522
                                                  30'd    5848    : data = 32'h    00835EB3    ;    //    srl x29 x6 x8      ====        srl t4, t1, s0
                                                  30'd    5849    : data = 32'h    397413B7    ;    //    lui x7 235329      ====        lui t2, 235329
                                                  30'd    5850    : data = 32'h    0111D313    ;    //    srli x6 x3 17      ====        srli t1, gp, 17
                                                  30'd    5851    : data = 32'h    40C38B33    ;    //    sub x22 x7 x12      ====        sub s6, t2, a2
                                                  30'd    5852    : data = 32'h    01E193B3    ;    //    sll x7 x3 x30      ====        sll t2, gp, t5
                                                  30'd    5853    : data = 32'h    FE4FF813    ;    //    andi x16 x31 -28      ====        andi a6, t6, -28
                                                  30'd    5854    : data = 32'h    3B50F713    ;    //    andi x14 x1 949      ====        andi a4, ra, 949
                                                  30'd    5855    : data = 32'h    0015F733    ;    //    and x14 x11 x1      ====        and a4, a1, ra
                                                  30'd    5856    : data = 32'h    C43BBE13    ;    //    sltiu x28 x23 -957      ====        sltiu t3, s7, -957
                                                  30'd    5857    : data = 32'h    3A4F19B7    ;    //    lui x19 238833      ====        lui s3, 238833
                                                  30'd    5858    : data = 32'h    93B53393    ;    //    sltiu x7 x10 -1733      ====        sltiu t2, a0, -1733
                                                  30'd    5859    : data = 32'h    012EE337    ;    //    lui x6 4846      ====        lui t1, 4846
                                                  30'd    5860    : data = 32'h    0008E193    ;    //    ori x3 x17 0      ====        ori gp, a7, 0
                                                  30'd    5861    : data = 32'h    008AF4B3    ;    //    and x9 x21 x8      ====        and s1, s5, s0
                                                  30'd    5862    : data = 32'h    4D9FCD17    ;    //    auipc x26 317948      ====        auipc s10, 317948
                                                  30'd    5863    : data = 32'h    41B65993    ;    //    srai x19 x12 27      ====        srai s3, a2, 27
                                                  30'd    5864    : data = 32'h    984E6C13    ;    //    ori x24 x28 -1660      ====        ori s8, t3, -1660
                                                  30'd    5865    : data = 32'h    0328AA17    ;    //    auipc x20 12938      ====        auipc s4, 12938
                                                  30'd    5866    : data = 32'h    013ADBB3    ;    //    srl x23 x21 x19      ====        srl s7, s5, s3
                                                  30'd    5867    : data = 32'h    40E80FB3    ;    //    sub x31 x16 x14      ====        sub t6, a6, a4
                                                  30'd    5868    : data = 32'h    00A69593    ;    //    slli x11 x13 10      ====        slli a1, a3, 10
                                                  30'd    5869    : data = 32'h    00412B33    ;    //    slt x22 x2 x4      ====        slt s6, sp, tp
                                                  30'd    5870    : data = 32'h    00C1C433    ;    //    xor x8 x3 x12      ====        xor s0, gp, a2
                                                  30'd    5871    : data = 32'h    D726ED93    ;    //    ori x27 x13 -654      ====        ori s11, a3, -654
                                                  30'd    5872    : data = 32'h    01769113    ;    //    slli x2 x13 23      ====        slli sp, a3, 23
                                                  30'd    5873    : data = 32'h    0F0E57B7    ;    //    lui x15 61669      ====        lui a5, 61669
                                                  30'd    5874    : data = 32'h    AE00BF93    ;    //    sltiu x31 x1 -1312      ====        sltiu t6, ra, -1312
                                                  30'd    5875    : data = 32'h    008ED333    ;    //    srl x6 x29 x8      ====        srl t1, t4, s0
                                                  30'd    5876    : data = 32'h    7991C393    ;    //    xori x7 x3 1945      ====        xori t2, gp, 1945
                                                  30'd    5877    : data = 32'h    B385A713    ;    //    slti x14 x11 -1224      ====        slti a4, a1, -1224
                                                  30'd    5878    : data = 32'h    EF8D4393    ;    //    xori x7 x26 -264      ====        xori t2, s10, -264
                                                  30'd    5879    : data = 32'h    2D683F93    ;    //    sltiu x31 x16 726      ====        sltiu t6, a6, 726
                                                  30'd    5880    : data = 32'h    F72B8613    ;    //    addi x12 x23 -142      ====        addi a2, s7, -142
                                                  30'd    5881    : data = 32'h    00AC0633    ;    //    add x12 x24 x10      ====        add a2, s8, a0
                                                  30'd    5882    : data = 32'h    018DC2B3    ;    //    xor x5 x27 x24      ====        xor t0, s11, s8
                                                  30'd    5883    : data = 32'h    6FC20093    ;    //    addi x1 x4 1788      ====        addi ra, tp, 1788
                                                  30'd    5884    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5885    : data = 32'h    01086AB3    ;    //    or x21 x16 x16      ====        or s5, a6, a6
                                                  30'd    5886    : data = 32'h    01F19613    ;    //    slli x12 x3 31      ====        slli a2, gp, 31
                                                  30'd    5887    : data = 32'h    BFF91D97    ;    //    auipc x27 786321      ====        auipc s11, 786321
                                                  30'd    5888    : data = 32'h    B0BCC613    ;    //    xori x12 x25 -1269      ====        xori a2, s9, -1269
                                                  30'd    5889    : data = 32'h    00438933    ;    //    add x18 x7 x4      ====        add s2, t2, tp
                                                  30'd    5890    : data = 32'h    00C145B3    ;    //    xor x11 x2 x12      ====        xor a1, sp, a2
                                                  30'd    5891    : data = 32'h    AF8E8B93    ;    //    addi x23 x29 -1288      ====        addi s7, t4, -1288
                                                  30'd    5892    : data = 32'h    009DC333    ;    //    xor x6 x27 x9      ====        xor t1, s11, s1
                                                  30'd    5893    : data = 32'h    7ED90A13    ;    //    addi x20 x18 2029      ====        addi s4, s2, 2029
                                                  30'd    5894    : data = 32'h    014A5AB3    ;    //    srl x21 x20 x20      ====        srl s5, s4, s4
                                                  30'd    5895    : data = 32'h    00425593    ;    //    srli x11 x4 4      ====        srli a1, tp, 4
                                                  30'd    5896    : data = 32'h    01845A93    ;    //    srli x21 x8 24      ====        srli s5, s0, 24
                                                  30'd    5897    : data = 32'h    013B2A33    ;    //    slt x20 x22 x19      ====        slt s4, s6, s3
                                                  30'd    5898    : data = 32'h    6E9301B7    ;    //    lui x3 452912      ====        lui gp, 452912
                                                  30'd    5899    : data = 32'h    408DD133    ;    //    sra x2 x27 x8      ====        sra sp, s11, s0
                                                  30'd    5900    : data = 32'h    44FC6313    ;    //    ori x6 x24 1103      ====        ori t1, s8, 1103
                                                  30'd    5901    : data = 32'h    415EED93    ;    //    ori x27 x29 1045      ====        ori s11, t4, 1045
                                                  30'd    5902    : data = 32'h    41565993    ;    //    srai x19 x12 21      ====        srai s3, a2, 21
                                                  30'd    5903    : data = 32'h    CFED0493    ;    //    addi x9 x26 -770      ====        addi s1, s10, -770
                                                  30'd    5904    : data = 32'h    00BC1713    ;    //    slli x14 x24 11      ====        slli a4, s8, 11
                                                  30'd    5905    : data = 32'h    0050FE33    ;    //    and x28 x1 x5      ====        and t3, ra, t0
                                                  30'd    5906    : data = 32'h    CF48BA13    ;    //    sltiu x20 x17 -780      ====        sltiu s4, a7, -780
                                                  30'd    5907    : data = 32'h    00C0EB33    ;    //    or x22 x1 x12      ====        or s6, ra, a2
                                                  30'd    5908    : data = 32'h    5ACA2093    ;    //    slti x1 x20 1452      ====        slti ra, s4, 1452
                                                  30'd    5909    : data = 32'h    01764333    ;    //    xor x6 x12 x23      ====        xor t1, a2, s7
                                                  30'd    5910    : data = 32'h    4073D9B3    ;    //    sra x19 x7 x7      ====        sra s3, t2, t2
                                                  30'd    5911    : data = 32'h    A51D7F97    ;    //    auipc x31 676311      ====        auipc t6, 676311
                                                  30'd    5912    : data = 32'h    00765C93    ;    //    srli x25 x12 7      ====        srli s9, a2, 7
                                                  30'd    5913    : data = 32'h    01231D93    ;    //    slli x27 x6 18      ====        slli s11, t1, 18
                                                  30'd    5914    : data = 32'h    95FEF713    ;    //    andi x14 x29 -1697      ====        andi a4, t4, -1697
                                                  30'd    5915    : data = 32'h    01489133    ;    //    sll x2 x17 x20      ====        sll sp, a7, s4
                                                  30'd    5916    : data = 32'h    0046C333    ;    //    xor x6 x13 x4      ====        xor t1, a3, tp
                                                  30'd    5917    : data = 32'h    34CE4D13    ;    //    xori x26 x28 844      ====        xori s10, t3, 844
                                                  30'd    5918    : data = 32'h    407F0633    ;    //    sub x12 x30 x7      ====        sub a2, t5, t2
                                                  30'd    5919    : data = 32'h    01C140B3    ;    //    xor x1 x2 x28      ====        xor ra, sp, t3
                                                  30'd    5920    : data = 32'h    0074B333    ;    //    sltu x6 x9 x7      ====        sltu t1, s1, t2
                                                  30'd    5921    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5922    : data = 32'h    01813733    ;    //    sltu x14 x2 x24      ====        sltu a4, sp, s8
                                                  30'd    5923    : data = 32'h    01F106B3    ;    //    add x13 x2 x31      ====        add a3, sp, t6
                                                  30'd    5924    : data = 32'h    00DCB633    ;    //    sltu x12 x25 x13      ====        sltu a2, s9, a3
                                                  30'd    5925    : data = 32'h    A7241CB7    ;    //    lui x25 684609      ====        lui s9, 684609
                                                  30'd    5926    : data = 32'h    018C9133    ;    //    sll x2 x25 x24      ====        sll sp, s9, s8
                                                  30'd    5927    : data = 32'h    D54C6793    ;    //    ori x15 x24 -684      ====        ori a5, s8, -684
                                                  30'd    5928    : data = 32'h    00D97DB3    ;    //    and x27 x18 x13      ====        and s11, s2, a3
                                                  30'd    5929    : data = 32'h    01AFDDB3    ;    //    srl x27 x31 x26      ====        srl s11, t6, s10
                                                  30'd    5930    : data = 32'h    00611E33    ;    //    sll x28 x2 x6      ====        sll t3, sp, t1
                                                  30'd    5931    : data = 32'h    D9808893    ;    //    addi x17 x1 -616      ====        addi a7, ra, -616
                                                  30'd    5932    : data = 32'h    41F45113    ;    //    srai x2 x8 31      ====        srai sp, s0, 31
                                                  30'd    5933    : data = 32'h    003576B3    ;    //    and x13 x10 x3      ====        and a3, a0, gp
                                                  30'd    5934    : data = 32'h    EB2F0813    ;    //    addi x16 x30 -334      ====        addi a6, t5, -334
                                                  30'd    5935    : data = 32'h    40D55D93    ;    //    srai x27 x10 13      ====        srai s11, a0, 13
                                                  30'd    5936    : data = 32'h    01E61033    ;    //    sll x0 x12 x30      ====        sll zero, a2, t5
                                                  30'd    5937    : data = 32'h    209BE4B7    ;    //    lui x9 133566      ====        lui s1, 133566
                                                  30'd    5938    : data = 32'h    00743133    ;    //    sltu x2 x8 x7      ====        sltu sp, s0, t2
                                                  30'd    5939    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5940    : data = 32'h    0051ECB3    ;    //    or x25 x3 x5      ====        or s9, gp, t0
                                                  30'd    5941    : data = 32'h    1917E713    ;    //    ori x14 x15 401      ====        ori a4, a5, 401
                                                  30'd    5942    : data = 32'h    9EA0EC93    ;    //    ori x25 x1 -1558      ====        ori s9, ra, -1558
                                                  30'd    5943    : data = 32'h    01EC5493    ;    //    srli x9 x24 30      ====        srli s1, s8, 30
                                                  30'd    5944    : data = 32'h    0114D4B3    ;    //    srl x9 x9 x17      ====        srl s1, s1, a7
                                                  30'd    5945    : data = 32'h    F6242893    ;    //    slti x17 x8 -158      ====        slti a7, s0, -158
                                                  30'd    5946    : data = 32'h    C27CB113    ;    //    sltiu x2 x25 -985      ====        sltiu sp, s9, -985
                                                  30'd    5947    : data = 32'h    E20C0693    ;    //    addi x13 x24 -480      ====        addi a3, s8, -480
                                                  30'd    5948    : data = 32'h    01F11433    ;    //    sll x8 x2 x31      ====        sll s0, sp, t6
                                                  30'd    5949    : data = 32'h    01E95813    ;    //    srli x16 x18 30      ====        srli a6, s2, 30
                                                  30'd    5950    : data = 32'h    F86FA093    ;    //    slti x1 x31 -122      ====        slti ra, t6, -122
                                                  30'd    5951    : data = 32'h    001D52B3    ;    //    srl x5 x26 x1      ====        srl t0, s10, ra
                                                  30'd    5952    : data = 32'h    0025B4B3    ;    //    sltu x9 x11 x2      ====        sltu s1, a1, sp
                                                  30'd    5953    : data = 32'h    404A5D93    ;    //    srai x27 x20 4      ====        srai s11, s4, 4
                                                  30'd    5954    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5955    : data = 32'h    774CC393    ;    //    xori x7 x25 1908      ====        xori t2, s9, 1908
                                                  30'd    5956    : data = 32'h    41800A33    ;    //    sub x20 x0 x24      ====        sub s4, zero, s8
                                                  30'd    5957    : data = 32'h    419C8EB3    ;    //    sub x29 x25 x25      ====        sub t4, s9, s9
                                                  30'd    5958    : data = 32'h    7341CC17    ;    //    auipc x24 472092      ====        auipc s8, 472092
                                                  30'd    5959    : data = 32'h    416255B3    ;    //    sra x11 x4 x22      ====        sra a1, tp, s6
                                                  30'd    5960    : data = 32'h    00F51D13    ;    //    slli x26 x10 15      ====        slli s10, a0, 15
                                                  30'd    5961    : data = 32'h    00F2EA33    ;    //    or x20 x5 x15      ====        or s4, t0, a5
                                                  30'd    5962    : data = 32'h    402F5C13    ;    //    srai x24 x30 2      ====        srai s8, t5, 2
                                                  30'd    5963    : data = 32'h    0076E733    ;    //    or x14 x13 x7      ====        or a4, a3, t2
                                                  30'd    5964    : data = 32'h    001CFEB3    ;    //    and x29 x25 x1      ====        and t4, s9, ra
                                                  30'd    5965    : data = 32'h    403A87B3    ;    //    sub x15 x21 x3      ====        sub a5, s5, gp
                                                  30'd    5966    : data = 32'h    05BF1B17    ;    //    auipc x22 23537      ====        auipc s6, 23537
                                                  30'd    5967    : data = 32'h    40A404B3    ;    //    sub x9 x8 x10      ====        sub s1, s0, a0
                                                  30'd    5968    : data = 32'h    0100F9B3    ;    //    and x19 x1 x16      ====        and s3, ra, a6
                                                  30'd    5969    : data = 32'h    C6674913    ;    //    xori x18 x14 -922      ====        xori s2, a4, -922
                                                  30'd    5970    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5971    : data = 32'h    017E1133    ;    //    sll x2 x28 x23      ====        sll sp, t3, s7
                                                  30'd    5972    : data = 32'h    D7B94293    ;    //    xori x5 x18 -645      ====        xori t0, s2, -645
                                                  30'd    5973    : data = 32'h    01F9F733    ;    //    and x14 x19 x31      ====        and a4, s3, t6
                                                  30'd    5974    : data = 32'h    00F4B633    ;    //    sltu x12 x9 x15      ====        sltu a2, s1, a5
                                                  30'd    5975    : data = 32'h    41C75813    ;    //    srai x16 x14 28      ====        srai a6, a4, 28
                                                  30'd    5976    : data = 32'h    01021F93    ;    //    slli x31 x4 16      ====        slli t6, tp, 16
                                                  30'd    5977    : data = 32'h    063CAC13    ;    //    slti x24 x25 99      ====        slti s8, s9, 99
                                                  30'd    5978    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5979    : data = 32'h    03ED4593    ;    //    xori x11 x26 62      ====        xori a1, s10, 62
                                                  30'd    5980    : data = 32'h    6F90E493    ;    //    ori x9 x1 1785      ====        ori s1, ra, 1785
                                                  30'd    5981    : data = 32'h    9D2DAD93    ;    //    slti x27 x27 -1582      ====        slti s11, s11, -1582
                                                  30'd    5982    : data = 32'h    7BB0E193    ;    //    ori x3 x1 1979      ====        ori gp, ra, 1979
                                                  30'd    5983    : data = 32'h    5A008C13    ;    //    addi x24 x1 1440      ====        addi s8, ra, 1440
                                                  30'd    5984    : data = 32'h    40B65713    ;    //    srai x14 x12 11      ====        srai a4, a2, 11
                                                  30'd    5985    : data = 32'h    3ACEED13    ;    //    ori x26 x29 940      ====        ori s10, t4, 940
                                                  30'd    5986    : data = 32'h    002F28B3    ;    //    slt x17 x30 x2      ====        slt a7, t5, sp
                                                  30'd    5987    : data = 32'h    7985F397    ;    //    auipc x7 497759      ====        auipc t2, 497759
                                                  30'd    5988    : data = 32'h    01E99C93    ;    //    slli x25 x19 30      ====        slli s9, s3, 30
                                                  30'd    5989    : data = 32'h    01F33433    ;    //    sltu x8 x6 x31      ====        sltu s0, t1, t6
                                                  30'd    5990    : data = 32'h    9C752413    ;    //    slti x8 x10 -1593      ====        slti s0, a0, -1593
                                                  30'd    5991    : data = 32'h    01E096B3    ;    //    sll x13 x1 x30      ====        sll a3, ra, t5
                                                  30'd    5992    : data = 32'h    E91622B7    ;    //    lui x5 954722      ====        lui t0, 954722
                                                  30'd    5993    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5994    : data = 32'h    00A9CAB3    ;    //    xor x21 x19 x10      ====        xor s5, s3, a0
                                                  30'd    5995    : data = 32'h    01D0DA13    ;    //    srli x20 x1 29      ====        srli s4, ra, 29
                                                  30'd    5996    : data = 32'h    3BE72E17    ;    //    auipc x28 245362      ====        auipc t3, 245362
                                                  30'd    5997    : data = 32'h    CBE9F897    ;    //    auipc x17 835231      ====        auipc a7, 835231
                                                  30'd    5998    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    5999    : data = 32'h    BE8B1497    ;    //    auipc x9 780465      ====        auipc s1, 780465
                                                  30'd    6000    : data = 32'h    01043FB3    ;    //    sltu x31 x8 x16      ====        sltu t6, s0, a6
                                                  30'd    6001    : data = 32'h    412C5713    ;    //    srai x14 x24 18      ====        srai a4, s8, 18
                                                  30'd    6002    : data = 32'h    013061B3    ;    //    or x3 x0 x19      ====        or gp, zero, s3
                                                  30'd    6003    : data = 32'h    690E6C93    ;    //    ori x25 x28 1680      ====        ori s9, t3, 1680
                                                  30'd    6004    : data = 32'h    0DC10C13    ;    //    addi x24 x2 220      ====        addi s8, sp, 220
                                                  30'd    6005    : data = 32'h    8BD8CE93    ;    //    xori x29 x17 -1859      ====        xori t4, a7, -1859
                                                  30'd    6006    : data = 32'h    014247B3    ;    //    xor x15 x4 x20      ====        xor a5, tp, s4
                                                  30'd    6007    : data = 32'h    4005D733    ;    //    sra x14 x11 x0      ====        sra a4, a1, zero
                                                  30'd    6008    : data = 32'h    00CF4AB3    ;    //    xor x21 x30 x12      ====        xor s5, t5, a2
                                                  30'd    6009    : data = 32'h    F7EE1F97    ;    //    auipc x31 1015521      ====        auipc t6, 1015521
                                                  30'd    6010    : data = 32'h    003FDD93    ;    //    srli x27 x31 3      ====        srli s11, t6, 3
                                                  30'd    6011    : data = 32'h    006612B3    ;    //    sll x5 x12 x6      ====        sll t0, a2, t1
                                                  30'd    6012    : data = 32'h    40A7D493    ;    //    srai x9 x15 10      ====        srai s1, a5, 10
                                                  30'd    6013    : data = 32'h    002C9A13    ;    //    slli x20 x25 2      ====        slli s4, s9, 2
                                                  30'd    6014    : data = 32'h    001C6AB3    ;    //    or x21 x24 x1      ====        or s5, s8, ra
                                                  30'd    6015    : data = 32'h    0154B2B3    ;    //    sltu x5 x9 x21      ====        sltu t0, s1, s5
                                                  30'd    6016    : data = 32'h    334D0813    ;    //    addi x16 x26 820      ====        addi a6, s10, 820
                                                  30'd    6017    : data = 32'h    40BAD3B3    ;    //    sra x7 x21 x11      ====        sra t2, s5, a1
                                                  30'd    6018    : data = 32'h    66A04713    ;    //    xori x14 x0 1642      ====        xori a4, zero, 1642
                                                  30'd    6019    : data = 32'h    015CF433    ;    //    and x8 x25 x21      ====        and s0, s9, s5
                                                  30'd    6020    : data = 32'h    A14A8413    ;    //    addi x8 x21 -1516      ====        addi s0, s5, -1516
                                                  30'd    6021    : data = 32'h    00DA75B3    ;    //    and x11 x20 x13      ====        and a1, s4, a3
                                                  30'd    6022    : data = 32'h    00DC6733    ;    //    or x14 x24 x13      ====        or a4, s8, a3
                                                  30'd    6023    : data = 32'h    41265913    ;    //    srai x18 x12 18      ====        srai s2, a2, 18
                                                  30'd    6024    : data = 32'h    40A05393    ;    //    srai x7 x0 10      ====        srai t2, zero, 10
                                                  30'd    6025    : data = 32'h    8260F393    ;    //    andi x7 x1 -2010      ====        andi t2, ra, -2010
                                                  30'd    6026    : data = 32'h    00C6EEB3    ;    //    or x29 x13 x12      ====        or t4, a3, a2
                                                  30'd    6027    : data = 32'h    00969493    ;    //    slli x9 x13 9      ====        slli s1, a3, 9
                                                  30'd    6028    : data = 32'h    0169EC33    ;    //    or x24 x19 x22      ====        or s8, s3, s6
                                                  30'd    6029    : data = 32'h    40B783B3    ;    //    sub x7 x15 x11      ====        sub t2, a5, a1
                                                  30'd    6030    : data = 32'h    000768B3    ;    //    or x17 x14 x0      ====        or a7, a4, zero
                                                  30'd    6031    : data = 32'h    348FA613    ;    //    slti x12 x31 840      ====        slti a2, t6, 840
                                                  30'd    6032    : data = 32'h    01100C93    ;    //    addi x25 x0 17      ====        addi s9, zero, 17
                                                  30'd    6033    : data = 32'h    F245AC37    ;    //    lui x24 992346      ====        lui s8, 992346
                                                  30'd    6034    : data = 32'h    0CD24013    ;    //    xori x0 x4 205      ====        xori zero, tp, 205
                                                  30'd    6035    : data = 32'h    1D3F0D93    ;    //    addi x27 x30 467      ====        addi s11, t5, 467
                                                  30'd    6036    : data = 32'h    01805B13    ;    //    srli x22 x0 24      ====        srli s6, zero, 24
                                                  30'd    6037    : data = 32'h    015BD2B3    ;    //    srl x5 x23 x21      ====        srl t0, s7, s5
                                                  30'd    6038    : data = 32'h    000492B3    ;    //    sll x5 x9 x0      ====        sll t0, s1, zero
                                                  30'd    6039    : data = 32'h    1F35B793    ;    //    sltiu x15 x11 499      ====        sltiu a5, a1, 499
                                                  30'd    6040    : data = 32'h    01B7C1B3    ;    //    xor x3 x15 x27      ====        xor gp, a5, s11
                                                  30'd    6041    : data = 32'h    019E3633    ;    //    sltu x12 x28 x25      ====        sltu a2, t3, s9
                                                  30'd    6042    : data = 32'h    0090D5B3    ;    //    srl x11 x1 x9      ====        srl a1, ra, s1
                                                  30'd    6043    : data = 32'h    5E07C113    ;    //    xori x2 x15 1504      ====        xori sp, a5, 1504
                                                  30'd    6044    : data = 32'h    01F719B3    ;    //    sll x19 x14 x31      ====        sll s3, a4, t6
                                                  30'd    6045    : data = 32'h    01F1DDB3    ;    //    srl x27 x3 x31      ====        srl s11, gp, t6
                                                  30'd    6046    : data = 32'h    9BC5C713    ;    //    xori x14 x11 -1604      ====        xori a4, a1, -1604
                                                  30'd    6047    : data = 32'h    23CB2093    ;    //    slti x1 x22 572      ====        slti ra, s6, 572
                                                  30'd    6048    : data = 32'h    7FC34893    ;    //    xori x17 x6 2044      ====        xori a7, t1, 2044
                                                  30'd    6049    : data = 32'h    00F29793    ;    //    slli x15 x5 15      ====        slli a5, t0, 15
                                                  30'd    6050    : data = 32'h    CDF78B13    ;    //    addi x22 x15 -801      ====        addi s6, a5, -801
                                                  30'd    6051    : data = 32'h    541D8E13    ;    //    addi x28 x27 1345      ====        addi t3, s11, 1345
                                                  30'd    6052    : data = 32'h    0162D9B3    ;    //    srl x19 x5 x22      ====        srl s3, t0, s6
                                                  30'd    6053    : data = 32'h    405E5913    ;    //    srai x18 x28 5      ====        srai s2, t3, 5
                                                  30'd    6054    : data = 32'h    019F1BB3    ;    //    sll x23 x30 x25      ====        sll s7, t5, s9
                                                  30'd    6055    : data = 32'h    79B1E493    ;    //    ori x9 x3 1947      ====        ori s1, gp, 1947
                                                  30'd    6056    : data = 32'h    00A25633    ;    //    srl x12 x4 x10      ====        srl a2, tp, a0
                                                  30'd    6057    : data = 32'h    00E5CBB3    ;    //    xor x23 x11 x14      ====        xor s7, a1, a4
                                                  30'd    6058    : data = 32'h    410152B3    ;    //    sra x5 x2 x16      ====        sra t0, sp, a6
                                                  30'd    6059    : data = 32'h    01C25B33    ;    //    srl x22 x4 x28      ====        srl s6, tp, t3
                                                  30'd    6060    : data = 32'h    401C02B3    ;    //    sub x5 x24 x1      ====        sub t0, s8, ra
                                                  30'd    6061    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6062    : data = 32'h    414E0833    ;    //    sub x16 x28 x20      ====        sub a6, t3, s4
                                                  30'd    6063    : data = 32'h    00785A13    ;    //    srli x20 x16 7      ====        srli s4, a6, 7
                                                  30'd    6064    : data = 32'h    40205333    ;    //    sra x6 x0 x2      ====        sra t1, zero, sp
                                                  30'd    6065    : data = 32'h    6A7F62B7    ;    //    lui x5 436214      ====        lui t0, 436214
                                                  30'd    6066    : data = 32'h    0A1AF793    ;    //    andi x15 x21 161      ====        andi a5, s5, 161
                                                  30'd    6067    : data = 32'h    8A7E8593    ;    //    addi x11 x29 -1881      ====        addi a1, t4, -1881
                                                  30'd    6068    : data = 32'h    415D0033    ;    //    sub x0 x26 x21      ====        sub zero, s10, s5
                                                  30'd    6069    : data = 32'h    00A610B3    ;    //    sll x1 x12 x10      ====        sll ra, a2, a0
                                                  30'd    6070    : data = 32'h    78FB7093    ;    //    andi x1 x22 1935      ====        andi ra, s6, 1935
                                                  30'd    6071    : data = 32'h    01469593    ;    //    slli x11 x13 20      ====        slli a1, a3, 20
                                                  30'd    6072    : data = 32'h    30878593    ;    //    addi x11 x15 776      ====        addi a1, a5, 776
                                                  30'd    6073    : data = 32'h    D47A6C93    ;    //    ori x25 x20 -697      ====        ori s9, s4, -697
                                                  30'd    6074    : data = 32'h    0044FE33    ;    //    and x28 x9 x4      ====        and t3, s1, tp
                                                  30'd    6075    : data = 32'h    010B5F93    ;    //    srli x31 x22 16      ====        srli t6, s6, 16
                                                  30'd    6076    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6077    : data = 32'h    A5197593    ;    //    andi x11 x18 -1455      ====        andi a1, s2, -1455
                                                  30'd    6078    : data = 32'h    00959613    ;    //    slli x12 x11 9      ====        slli a2, a1, 9
                                                  30'd    6079    : data = 32'h    00259B13    ;    //    slli x22 x11 2      ====        slli s6, a1, 2
                                                  30'd    6080    : data = 32'h    00AEABB3    ;    //    slt x23 x29 x10      ====        slt s7, t4, a0
                                                  30'd    6081    : data = 32'h    C894F813    ;    //    andi x16 x9 -887      ====        andi a6, s1, -887
                                                  30'd    6082    : data = 32'h    002ED9B3    ;    //    srl x19 x29 x2      ====        srl s3, t4, sp
                                                  30'd    6083    : data = 32'h    8CDCAE93    ;    //    slti x29 x25 -1843      ====        slti t4, s9, -1843
                                                  30'd    6084    : data = 32'h    00D421B3    ;    //    slt x3 x8 x13      ====        slt gp, s0, a3
                                                  30'd    6085    : data = 32'h    000F9893    ;    //    slli x17 x31 0      ====        slli a7, t6, 0
                                                  30'd    6086    : data = 32'h    00A017B3    ;    //    sll x15 x0 x10      ====        sll a5, zero, a0
                                                  30'd    6087    : data = 32'h    002E78B3    ;    //    and x17 x28 x2      ====        and a7, t3, sp
                                                  30'd    6088    : data = 32'h    418151B3    ;    //    sra x3 x2 x24      ====        sra gp, sp, s8
                                                  30'd    6089    : data = 32'h    413188B3    ;    //    sub x17 x3 x19      ====        sub a7, gp, s3
                                                  30'd    6090    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6091    : data = 32'h    01F2D793    ;    //    srli x15 x5 31      ====        srli a5, t0, 31
                                                  30'd    6092    : data = 32'h    011B1FB3    ;    //    sll x31 x22 x17      ====        sll t6, s6, a7
                                                  30'd    6093    : data = 32'h    003065B3    ;    //    or x11 x0 x3      ====        or a1, zero, gp
                                                  30'd    6094    : data = 32'h    94FE4E93    ;    //    xori x29 x28 -1713      ====        xori t4, t3, -1713
                                                  30'd    6095    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6096    : data = 32'h    00E10033    ;    //    add x0 x2 x14      ====        add zero, sp, a4
                                                  30'd    6097    : data = 32'h    007DB733    ;    //    sltu x14 x27 x7      ====        sltu a4, s11, t2
                                                  30'd    6098    : data = 32'h    00268FB3    ;    //    add x31 x13 x2      ====        add t6, a3, sp
                                                  30'd    6099    : data = 32'h    CA5FBD93    ;    //    sltiu x27 x31 -859      ====        sltiu s11, t6, -859
                                                  30'd    6100    : data = 32'h    00A599B3    ;    //    sll x19 x11 x10      ====        sll s3, a1, a0
                                                  30'd    6101    : data = 32'h    01EA7133    ;    //    and x2 x20 x30      ====        and sp, s4, t5
                                                  30'd    6102    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6103    : data = 32'h    402B84B3    ;    //    sub x9 x23 x2      ====        sub s1, s7, sp
                                                  30'd    6104    : data = 32'h    5A768813    ;    //    addi x16 x13 1447      ====        addi a6, a3, 1447
                                                  30'd    6105    : data = 32'h    41638DB3    ;    //    sub x27 x7 x22      ====        sub s11, t2, s6
                                                  30'd    6106    : data = 32'h    01F134B3    ;    //    sltu x9 x2 x31      ====        sltu s1, sp, t6
                                                  30'd    6107    : data = 32'h    C9B2B593    ;    //    sltiu x11 x5 -869      ====        sltiu a1, t0, -869
                                                  30'd    6108    : data = 32'h    00E78EB3    ;    //    add x29 x15 x14      ====        add t4, a5, a4
                                                  30'd    6109    : data = 32'h    404DDB93    ;    //    srai x23 x27 4      ====        srai s7, s11, 4
                                                  30'd    6110    : data = 32'h    018E0733    ;    //    add x14 x28 x24      ====        add a4, t3, s8
                                                  30'd    6111    : data = 32'h    00F37933    ;    //    and x18 x6 x15      ====        and s2, t1, a5
                                                  30'd    6112    : data = 32'h    B4328E13    ;    //    addi x28 x5 -1213      ====        addi t3, t0, -1213
                                                  30'd    6113    : data = 32'h    01677E33    ;    //    and x28 x14 x22      ====        and t3, a4, s6
                                                  30'd    6114    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6115    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6116    : data = 32'h    196D2893    ;    //    slti x17 x26 406      ====        slti a7, s10, 406
                                                  30'd    6117    : data = 32'h    011AE4B3    ;    //    or x9 x21 x17      ====        or s1, s5, a7
                                                  30'd    6118    : data = 32'h    01A97EB3    ;    //    and x29 x18 x26      ====        and t4, s2, s10
                                                  30'd    6119    : data = 32'h    66D8CE93    ;    //    xori x29 x17 1645      ====        xori t4, a7, 1645
                                                  30'd    6120    : data = 32'h    003DDCB3    ;    //    srl x25 x27 x3      ====        srl s9, s11, gp
                                                  30'd    6121    : data = 32'h    00239813    ;    //    slli x16 x7 2      ====        slli a6, t2, 2
                                                  30'd    6122    : data = 32'h    005D5013    ;    //    srli x0 x26 5      ====        srli zero, s10, 5
                                                  30'd    6123    : data = 32'h    00ABD893    ;    //    srli x17 x23 10      ====        srli a7, s7, 10
                                                  30'd    6124    : data = 32'h    013B3C33    ;    //    sltu x24 x22 x19      ====        sltu s8, s6, s3
                                                  30'd    6125    : data = 32'h    0175ACB3    ;    //    slt x25 x11 x23      ====        slt s9, a1, s7
                                                  30'd    6126    : data = 32'h    9CAB8493    ;    //    addi x9 x23 -1590      ====        addi s1, s7, -1590
                                                  30'd    6127    : data = 32'h    003C4E33    ;    //    xor x28 x24 x3      ====        xor t3, s8, gp
                                                  30'd    6128    : data = 32'h    00180133    ;    //    add x2 x16 x1      ====        add sp, a6, ra
                                                  30'd    6129    : data = 32'h    40DD5693    ;    //    srai x13 x26 13      ====        srai a3, s10, 13
                                                  30'd    6130    : data = 32'h    0116B8B3    ;    //    sltu x17 x13 x17      ====        sltu a7, a3, a7
                                                  30'd    6131    : data = 32'h    49166793    ;    //    ori x15 x12 1169      ====        ori a5, a2, 1169
                                                  30'd    6132    : data = 32'h    00B6C033    ;    //    xor x0 x13 x11      ====        xor zero, a3, a1
                                                  30'd    6133    : data = 32'h    EF4A6713    ;    //    ori x14 x20 -268      ====        ori a4, s4, -268
                                                  30'd    6134    : data = 32'h    01381113    ;    //    slli x2 x16 19      ====        slli sp, a6, 19
                                                  30'd    6135    : data = 32'h    F374E993    ;    //    ori x19 x9 -201      ====        ori s3, s1, -201
                                                  30'd    6136    : data = 32'h    35038613    ;    //    addi x12 x7 848      ====        addi a2, t2, 848
                                                  30'd    6137    : data = 32'h    00E31C93    ;    //    slli x25 x6 14      ====        slli s9, t1, 14
                                                  30'd    6138    : data = 32'h    407B5B13    ;    //    srai x22 x22 7      ====        srai s6, s6, 7
                                                  30'd    6139    : data = 32'h    00601633    ;    //    sll x12 x0 x6      ====        sll a2, zero, t1
                                                  30'd    6140    : data = 32'h    794F5317    ;    //    auipc x6 496885      ====        auipc t1, 496885
                                                  30'd    6141    : data = 32'h    01C6F0B3    ;    //    and x1 x13 x28      ====        and ra, a3, t3
                                                  30'd    6142    : data = 32'h    39CA7293    ;    //    andi x5 x20 924      ====        andi t0, s4, 924
                                                  30'd    6143    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6144    : data = 32'h    40530D33    ;    //    sub x26 x6 x5      ====        sub s10, t1, t0
                                                  30'd    6145    : data = 32'h    008B6733    ;    //    or x14 x22 x8      ====        or a4, s6, s0
                                                  30'd    6146    : data = 32'h    487FCF93    ;    //    xori x31 x31 1159      ====        xori t6, t6, 1159
                                                  30'd    6147    : data = 32'h    01491193    ;    //    slli x3 x18 20      ====        slli gp, s2, 20
                                                  30'd    6148    : data = 32'h    00709E33    ;    //    sll x28 x1 x7      ====        sll t3, ra, t2
                                                  30'd    6149    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6150    : data = 32'h    003A5913    ;    //    srli x18 x20 3      ====        srli s2, s4, 3
                                                  30'd    6151    : data = 32'h    D7387317    ;    //    auipc x6 881543      ====        auipc t1, 881543
                                                  30'd    6152    : data = 32'h    018E5813    ;    //    srli x16 x28 24      ====        srli a6, t3, 24
                                                  30'd    6153    : data = 32'h    00DD6833    ;    //    or x16 x26 x13      ====        or a6, s10, a3
                                                  30'd    6154    : data = 32'h    F396C713    ;    //    xori x14 x13 -199      ====        xori a4, a3, -199
                                                  30'd    6155    : data = 32'h    D582C913    ;    //    xori x18 x5 -680      ====        xori s2, t0, -680
                                                  30'd    6156    : data = 32'h    95D2F317    ;    //    auipc x6 613679      ====        auipc t1, 613679
                                                  30'd    6157    : data = 32'h    EA2D3C17    ;    //    auipc x24 959187      ====        auipc s8, 959187
                                                  30'd    6158    : data = 32'h    01D7E5B3    ;    //    or x11 x15 x29      ====        or a1, a5, t4
                                                  30'd    6159    : data = 32'h    21F89C17    ;    //    auipc x24 139145      ====        auipc s8, 139145
                                                  30'd    6160    : data = 32'h    E6917EB7    ;    //    lui x29 944407      ====        lui t4, 944407
                                                  30'd    6161    : data = 32'h    008F5E33    ;    //    srl x28 x30 x8      ====        srl t3, t5, s0
                                                  30'd    6162    : data = 32'h    4054DB93    ;    //    srai x23 x9 5      ====        srai s7, s1, 5
                                                  30'd    6163    : data = 32'h    0153C733    ;    //    xor x14 x7 x21      ====        xor a4, t2, s5
                                                  30'd    6164    : data = 32'h    00780AB3    ;    //    add x21 x16 x7      ====        add s5, a6, t2
                                                  30'd    6165    : data = 32'h    00DC9FB3    ;    //    sll x31 x25 x13      ====        sll t6, s9, a3
                                                  30'd    6166    : data = 32'h    012B88B3    ;    //    add x17 x23 x18      ====        add a7, s7, s2
                                                  30'd    6167    : data = 32'h    69464093    ;    //    xori x1 x12 1684      ====        xori ra, a2, 1684
                                                  30'd    6168    : data = 32'h    007994B3    ;    //    sll x9 x19 x7      ====        sll s1, s3, t2
                                                  30'd    6169    : data = 32'h    40A6DE13    ;    //    srai x28 x13 10      ====        srai t3, a3, 10
                                                  30'd    6170    : data = 32'h    CF7C2B13    ;    //    slti x22 x24 -777      ====        slti s6, s8, -777
                                                  30'd    6171    : data = 32'h    009CA5B3    ;    //    slt x11 x25 x9      ====        slt a1, s9, s1
                                                  30'd    6172    : data = 32'h    00C45733    ;    //    srl x14 x8 x12      ====        srl a4, s0, a2
                                                  30'd    6173    : data = 32'h    DD677293    ;    //    andi x5 x14 -554      ====        andi t0, a4, -554
                                                  30'd    6174    : data = 32'h    002EDE13    ;    //    srli x28 x29 2      ====        srli t3, t4, 2
                                                  30'd    6175    : data = 32'h    005CF8B3    ;    //    and x17 x25 x5      ====        and a7, s9, t0
                                                  30'd    6176    : data = 32'h    78630313    ;    //    addi x6 x6 1926      ====        addi t1, t1, 1926
                                                  30'd    6177    : data = 32'h    01B27A33    ;    //    and x20 x4 x27      ====        and s4, tp, s11
                                                  30'd    6178    : data = 32'h    EA622097    ;    //    auipc x1 960034      ====        auipc ra, 960034
                                                  30'd    6179    : data = 32'h    3A614C13    ;    //    xori x24 x2 934      ====        xori s8, sp, 934
                                                  30'd    6180    : data = 32'h    0183A033    ;    //    slt x0 x7 x24      ====        slt zero, t2, s8
                                                  30'd    6181    : data = 32'h    ABFC6613    ;    //    ori x12 x24 -1345      ====        ori a2, s8, -1345
                                                  30'd    6182    : data = 32'h    00AADF93    ;    //    srli x31 x21 10      ====        srli t6, s5, 10
                                                  30'd    6183    : data = 32'h    DB343C97    ;    //    auipc x25 897859      ====        auipc s9, 897859
                                                  30'd    6184    : data = 32'h    E69FBC93    ;    //    sltiu x25 x31 -407      ====        sltiu s9, t6, -407
                                                  30'd    6185    : data = 32'h    1D0B8A13    ;    //    addi x20 x23 464      ====        addi s4, s7, 464
                                                  30'd    6186    : data = 32'h    00A7D113    ;    //    srli x2 x15 10      ====        srli sp, a5, 10
                                                  30'd    6187    : data = 32'h    CBD63B93    ;    //    sltiu x23 x12 -835      ====        sltiu s7, a2, -835
                                                  30'd    6188    : data = 32'h    41885793    ;    //    srai x15 x16 24      ====        srai a5, a6, 24
                                                  30'd    6189    : data = 32'h    005F2933    ;    //    slt x18 x30 x5      ====        slt s2, t5, t0
                                                  30'd    6190    : data = 32'h    01823333    ;    //    sltu x6 x4 x24      ====        sltu t1, tp, s8
                                                  30'd    6191    : data = 32'h    E52B8893    ;    //    addi x17 x23 -430      ====        addi a7, s7, -430
                                                  30'd    6192    : data = 32'h    01C5C833    ;    //    xor x16 x11 x28      ====        xor a6, a1, t3
                                                  30'd    6193    : data = 32'h    68686313    ;    //    ori x6 x16 1670      ====        ori t1, a6, 1670
                                                  30'd    6194    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6195    : data = 32'h    00FC6BB3    ;    //    or x23 x24 x15      ====        or s7, s8, a5
                                                  30'd    6196    : data = 32'h    610CE893    ;    //    ori x17 x25 1552      ====        ori a7, s9, 1552
                                                  30'd    6197    : data = 32'h    0145AAB3    ;    //    slt x21 x11 x20      ====        slt s5, a1, s4
                                                  30'd    6198    : data = 32'h    01915013    ;    //    srli x0 x2 25      ====        srli zero, sp, 25
                                                  30'd    6199    : data = 32'h    0006D613    ;    //    srli x12 x13 0      ====        srli a2, a3, 0
                                                  30'd    6200    : data = 32'h    0D47F813    ;    //    andi x16 x15 212      ====        andi a6, a5, 212
                                                  30'd    6201    : data = 32'h    0110E1B3    ;    //    or x3 x1 x17      ====        or gp, ra, a7
                                                  30'd    6202    : data = 32'h    018531B3    ;    //    sltu x3 x10 x24      ====        sltu gp, a0, s8
                                                  30'd    6203    : data = 32'h    4143DC33    ;    //    sra x24 x7 x20      ====        sra s8, t2, s4
                                                  30'd    6204    : data = 32'h    41A3D6B3    ;    //    sra x13 x7 x26      ====        sra a3, t2, s10
                                                  30'd    6205    : data = 32'h    00D81193    ;    //    slli x3 x16 13      ====        slli gp, a6, 13
                                                  30'd    6206    : data = 32'h    41628433    ;    //    sub x8 x5 x22      ====        sub s0, t0, s6
                                                  30'd    6207    : data = 32'h    8E3F8097    ;    //    auipc x1 582648      ====        auipc ra, 582648
                                                  30'd    6208    : data = 32'h    0106FFB3    ;    //    and x31 x13 x16      ====        and t6, a3, a6
                                                  30'd    6209    : data = 32'h    B964A413    ;    //    slti x8 x9 -1130      ====        slti s0, s1, -1130
                                                  30'd    6210    : data = 32'h    4C524D93    ;    //    xori x27 x4 1221      ====        xori s11, tp, 1221
                                                  30'd    6211    : data = 32'h    D9D0CB93    ;    //    xori x23 x1 -611      ====        xori s7, ra, -611
                                                  30'd    6212    : data = 32'h    008D5593    ;    //    srli x11 x26 8      ====        srli a1, s10, 8
                                                  30'd    6213    : data = 32'h    00A40FB3    ;    //    add x31 x8 x10      ====        add t6, s0, a0
                                                  30'd    6214    : data = 32'h    0074CAB3    ;    //    xor x21 x9 x7      ====        xor s5, s1, t2
                                                  30'd    6215    : data = 32'h    06BA8693    ;    //    addi x13 x21 107      ====        addi a3, s5, 107
                                                  30'd    6216    : data = 32'h    8B7CBB13    ;    //    sltiu x22 x25 -1865      ====        sltiu s6, s9, -1865
                                                  30'd    6217    : data = 32'h    585C2813    ;    //    slti x16 x24 1413      ====        slti a6, s8, 1413
                                                  30'd    6218    : data = 32'h    00A0E5B3    ;    //    or x11 x1 x10      ====        or a1, ra, a0
                                                  30'd    6219    : data = 32'h    010910B3    ;    //    sll x1 x18 x16      ====        sll ra, s2, a6
                                                  30'd    6220    : data = 32'h    01430633    ;    //    add x12 x6 x20      ====        add a2, t1, s4
                                                  30'd    6221    : data = 32'h    01195293    ;    //    srli x5 x18 17      ====        srli t0, s2, 17
                                                  30'd    6222    : data = 32'h    00333033    ;    //    sltu x0 x6 x3      ====        sltu zero, t1, gp
                                                  30'd    6223    : data = 32'h    840DBE93    ;    //    sltiu x29 x27 -1984      ====        sltiu t4, s11, -1984
                                                  30'd    6224    : data = 32'h    01FE1413    ;    //    slli x8 x28 31      ====        slli s0, t3, 31
                                                  30'd    6225    : data = 32'h    001689B3    ;    //    add x19 x13 x1      ====        add s3, a3, ra
                                                  30'd    6226    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6227    : data = 32'h    01BF4133    ;    //    xor x2 x30 x27      ====        xor sp, t5, s11
                                                  30'd    6228    : data = 32'h    406D5733    ;    //    sra x14 x26 x6      ====        sra a4, s10, t1
                                                  30'd    6229    : data = 32'h    6192C593    ;    //    xori x11 x5 1561      ====        xori a1, t0, 1561
                                                  30'd    6230    : data = 32'h    417EDB13    ;    //    srai x22 x29 23      ====        srai s6, t4, 23
                                                  30'd    6231    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6232    : data = 32'h    81A6B413    ;    //    sltiu x8 x13 -2022      ====        sltiu s0, a3, -2022
                                                  30'd    6233    : data = 32'h    9F6D3897    ;    //    auipc x17 653011      ====        auipc a7, 653011
                                                  30'd    6234    : data = 32'h    3E14E413    ;    //    ori x8 x9 993      ====        ori s0, s1, 993
                                                  30'd    6235    : data = 32'h    01D93BB3    ;    //    sltu x23 x18 x29      ====        sltu s7, s2, t4
                                                  30'd    6236    : data = 32'h    41045313    ;    //    srai x6 x8 16      ====        srai t1, s0, 16
                                                  30'd    6237    : data = 32'h    D996BF93    ;    //    sltiu x31 x13 -615      ====        sltiu t6, a3, -615
                                                  30'd    6238    : data = 32'h    009895B3    ;    //    sll x11 x17 x9      ====        sll a1, a7, s1
                                                  30'd    6239    : data = 32'h    01E55693    ;    //    srli x13 x10 30      ====        srli a3, a0, 30
                                                  30'd    6240    : data = 32'h    416DDD13    ;    //    srai x26 x27 22      ====        srai s10, s11, 22
                                                  30'd    6241    : data = 32'h    9ABF7D13    ;    //    andi x26 x30 -1621      ====        andi s10, t5, -1621
                                                  30'd    6242    : data = 32'h    C898E013    ;    //    ori x0 x17 -887      ====        ori zero, a7, -887
                                                  30'd    6243    : data = 32'h    01C3D913    ;    //    srli x18 x7 28      ====        srli s2, t2, 28
                                                  30'd    6244    : data = 32'h    633ABA37    ;    //    lui x20 406443      ====        lui s4, 406443
                                                  30'd    6245    : data = 32'h    D60D17B7    ;    //    lui x15 876753      ====        lui a5, 876753
                                                  30'd    6246    : data = 32'h    00955D13    ;    //    srli x26 x10 9      ====        srli s10, a0, 9
                                                  30'd    6247    : data = 32'h    0131D293    ;    //    srli x5 x3 19      ====        srli t0, gp, 19
                                                  30'd    6248    : data = 32'h    00D68CB3    ;    //    add x25 x13 x13      ====        add s9, a3, a3
                                                  30'd    6249    : data = 32'h    41098A33    ;    //    sub x20 x19 x16      ====        sub s4, s3, a6
                                                  30'd    6250    : data = 32'h    00999693    ;    //    slli x13 x19 9      ====        slli a3, s3, 9
                                                  30'd    6251    : data = 32'h    417B87B3    ;    //    sub x15 x23 x23      ====        sub a5, s7, s7
                                                  30'd    6252    : data = 32'h    FBB52C13    ;    //    slti x24 x10 -69      ====        slti s8, a0, -69
                                                  30'd    6253    : data = 32'h    00A3C633    ;    //    xor x12 x7 x10      ====        xor a2, t2, a0
                                                  30'd    6254    : data = 32'h    011624B3    ;    //    slt x9 x12 x17      ====        slt s1, a2, a7
                                                  30'd    6255    : data = 32'h    01AED713    ;    //    srli x14 x29 26      ====        srli a4, t4, 26
                                                  30'd    6256    : data = 32'h    00391FB3    ;    //    sll x31 x18 x3      ====        sll t6, s2, gp
                                                  30'd    6257    : data = 32'h    AB6C6A93    ;    //    ori x21 x24 -1354      ====        ori s5, s8, -1354
                                                  30'd    6258    : data = 32'h    4150D013    ;    //    srai x0 x1 21      ====        srai zero, ra, 21
                                                  30'd    6259    : data = 32'h    01239813    ;    //    slli x16 x7 18      ====        slli a6, t2, 18
                                                  30'd    6260    : data = 32'h    15F5FA37    ;    //    lui x20 89951      ====        lui s4, 89951
                                                  30'd    6261    : data = 32'h    00BC6CB3    ;    //    or x25 x24 x11      ====        or s9, s8, a1
                                                  30'd    6262    : data = 32'h    AFF8A293    ;    //    slti x5 x17 -1281      ====        slti t0, a7, -1281
                                                  30'd    6263    : data = 32'h    40E85E93    ;    //    srai x29 x16 14      ====        srai t4, a6, 14
                                                  30'd    6264    : data = 32'h    000F3EB3    ;    //    sltu x29 x30 x0      ====        sltu t4, t5, zero
                                                  30'd    6265    : data = 32'h    294A6593    ;    //    ori x11 x20 660      ====        ori a1, s4, 660
                                                  30'd    6266    : data = 32'h    0030D713    ;    //    srli x14 x1 3      ====        srli a4, ra, 3
                                                  30'd    6267    : data = 32'h    009F2C33    ;    //    slt x24 x30 x9      ====        slt s8, t5, s1
                                                  30'd    6268    : data = 32'h    01004033    ;    //    xor x0 x0 x16      ====        xor zero, zero, a6
                                                  30'd    6269    : data = 32'h    70C0F493    ;    //    andi x9 x1 1804      ====        andi s1, ra, 1804
                                                  30'd    6270    : data = 32'h    01D3B033    ;    //    sltu x0 x7 x29      ====        sltu zero, t2, t4
                                                  30'd    6271    : data = 32'h    00A45293    ;    //    srli x5 x8 10      ====        srli t0, s0, 10
                                                  30'd    6272    : data = 32'h    40EBDAB3    ;    //    sra x21 x23 x14      ====        sra s5, s7, a4
                                                  30'd    6273    : data = 32'h    800002B7    ;    //    lui x5 524288      ====        li t0, 0x80000000 #start riscv_int_numeric_corner_stream_14
                                                  30'd    6274    : data = 32'h    00028293    ;    //    addi x5 x5 0      ====        li t0, 0x80000000 #start riscv_int_numeric_corner_stream_14
                                                  30'd    6275    : data = 32'h    00000693    ;    //    addi x13 x0 0      ====        li a3, 0x0
                                                  30'd    6276    : data = 32'h    00000393    ;    //    addi x7 x0 0      ====        li t2, 0x0
                                                  30'd    6277    : data = 32'h    B3CAFAB7    ;    //    lui x21 736431      ====        li s5, 0xb3cae956
                                                  30'd    6278    : data = 32'h    956A8A93    ;    //    addi x21 x21 -1706      ====        li s5, 0xb3cae956
                                                  30'd    6279    : data = 32'h    80000BB7    ;    //    lui x23 524288      ====        li s7, 0x80000000
                                                  30'd    6280    : data = 32'h    000B8B93    ;    //    addi x23 x23 0      ====        li s7, 0x80000000
                                                  30'd    6281    : data = 32'h    80000637    ;    //    lui x12 524288      ====        li a2, 0x80000000
                                                  30'd    6282    : data = 32'h    00060613    ;    //    addi x12 x12 0      ====        li a2, 0x80000000
                                                  30'd    6283    : data = 32'h    80000137    ;    //    lui x2 524288      ====        li sp, 0x80000000
                                                  30'd    6284    : data = 32'h    00010113    ;    //    addi x2 x2 0      ====        li sp, 0x80000000
                                                  30'd    6285    : data = 32'h    FFF00C13    ;    //    addi x24 x0 -1      ====        li s8, 0xffffffff
                                                  30'd    6286    : data = 32'h    80000837    ;    //    lui x16 524288      ====        li a6, 0x80000000
                                                  30'd    6287    : data = 32'h    00080813    ;    //    addi x16 x16 0      ====        li a6, 0x80000000
                                                  30'd    6288    : data = 32'h    FFF00E93    ;    //    addi x29 x0 -1      ====        li t4, 0xffffffff
                                                  30'd    6289    : data = 32'h    39938813    ;    //    addi x16 x7 921      ====        addi a6, t2, 921
                                                  30'd    6290    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6291    : data = 32'h    407C0133    ;    //    sub x2 x24 x7      ====        sub sp, s8, t2
                                                  30'd    6292    : data = 32'h    01568AB3    ;    //    add x21 x13 x21      ====        add s5, a3, s5
                                                  30'd    6293    : data = 32'h    3B7E8113    ;    //    addi x2 x29 951      ====        addi sp, t4, 951
                                                  30'd    6294    : data = 32'h    7C898EB7    ;    //    lui x29 510104      ====        lui t4, 510104
                                                  30'd    6295    : data = 32'h    BBD832B7    ;    //    lui x5 769411      ====        lui t0, 769411
                                                  30'd    6296    : data = 32'h    41DB8633    ;    //    sub x12 x23 x29      ====        sub a2, s7, t4
                                                  30'd    6297    : data = 32'h    62568A93    ;    //    addi x21 x13 1573      ====        addi s5, a3, 1573
                                                  30'd    6298    : data = 32'h    6F3B8293    ;    //    addi x5 x23 1779      ====        addi t0, s7, 1779
                                                  30'd    6299    : data = 32'h    6D52B117    ;    //    auipc x2 447787      ====        auipc sp, 447787
                                                  30'd    6300    : data = 32'h    41880833    ;    //    sub x16 x16 x24      ====        sub a6, a6, s8
                                                  30'd    6301    : data = 32'h    578A6637    ;    //    lui x12 358566      ====        lui a2, 358566
                                                  30'd    6302    : data = 32'h    156E8613    ;    //    addi x12 x29 342      ====        addi a2, t4, 342
                                                  30'd    6303    : data = 32'h    40C80833    ;    //    sub x16 x16 x12      ====        sub a6, a6, a2
                                                  30'd    6304    : data = 32'h    C2AB4637    ;    //    lui x12 797364      ====        lui a2, 797364
                                                  30'd    6305    : data = 32'h    32857C17    ;    //    auipc x24 206935      ====        auipc s8, 206935
                                                  30'd    6306    : data = 32'h    6E91F397    ;    //    auipc x7 452895      ====        auipc t2, 452895
                                                  30'd    6307    : data = 32'h    015C0833    ;    //    add x16 x24 x21      ====        add a6, s8, s5
                                                  30'd    6308    : data = 32'h    4B928813    ;    //    addi x16 x5 1209      ====        addi a6, t0, 1209
                                                  30'd    6309    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6310    : data = 32'h    010B8BB3    ;    //    add x23 x23 x16      ====        add s7, s7, a6
                                                  30'd    6311    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6312    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6313    : data = 32'h    017E8633    ;    //    add x12 x29 x23      ====        add a2, t4, s7
                                                  30'd    6314    : data = 32'h    3D84AC17    ;    //    auipc x24 251978      ====        auipc s8, 251978
                                                  30'd    6315    : data = 32'h    E93B8293    ;    //    addi x5 x23 -365      ====        addi t0, s7, -365
                                                  30'd    6316    : data = 32'h    438050EF    ;    //    jal x1 21560      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_14
                                                  30'd    6317    : data = 32'h    88892393    ;    //    slti x7 x18 -1912      ====        slti t2, s2, -1912
                                                  30'd    6318    : data = 32'h    01F778B3    ;    //    and x17 x14 x31      ====        and a7, a4, t6
                                                  30'd    6319    : data = 32'h    50DC0013    ;    //    addi x0 x24 1293      ====        addi zero, s8, 1293
                                                  30'd    6320    : data = 32'h    2516CDB7    ;    //    lui x27 151916      ====        lui s11, 151916
                                                  30'd    6321    : data = 32'h    0018C833    ;    //    xor x16 x17 x1      ====        xor a6, a7, ra
                                                  30'd    6322    : data = 32'h    01405593    ;    //    srli x11 x0 20      ====        srli a1, zero, 20
                                                  30'd    6323    : data = 32'h    41AD8033    ;    //    sub x0 x27 x26      ====        sub zero, s11, s10
                                                  30'd    6324    : data = 32'h    01B92833    ;    //    slt x16 x18 x27      ====        slt a6, s2, s11
                                                  30'd    6325    : data = 32'h    28192493    ;    //    slti x9 x18 641      ====        slti s1, s2, 641
                                                  30'd    6326    : data = 32'h    0320E693    ;    //    ori x13 x1 50      ====        ori a3, ra, 50
                                                  30'd    6327    : data = 32'h    00CAB5B3    ;    //    sltu x11 x21 x12      ====        sltu a1, s5, a2
                                                  30'd    6328    : data = 32'h    3B7980B7    ;    //    lui x1 243608      ====        lui ra, 243608
                                                  30'd    6329    : data = 32'h    2C1A3917    ;    //    auipc x18 180643      ====        auipc s2, 180643
                                                  30'd    6330    : data = 32'h    00764733    ;    //    xor x14 x12 x7      ====        xor a4, a2, t2
                                                  30'd    6331    : data = 32'h    09258E93    ;    //    addi x29 x11 146      ====        addi t4, a1, 146
                                                  30'd    6332    : data = 32'h    7F9C4993    ;    //    xori x19 x24 2041      ====        xori s3, s8, 2041
                                                  30'd    6333    : data = 32'h    E7BC2B13    ;    //    slti x22 x24 -389      ====        slti s6, s8, -389
                                                  30'd    6334    : data = 32'h    417DD313    ;    //    srai x6 x27 23      ====        srai t1, s11, 23
                                                  30'd    6335    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6336    : data = 32'h    246D6D13    ;    //    ori x26 x26 582      ====        ori s10, s10, 582
                                                  30'd    6337    : data = 32'h    01DAD5B3    ;    //    srl x11 x21 x29      ====        srl a1, s5, t4
                                                  30'd    6338    : data = 32'h    41780CB3    ;    //    sub x25 x16 x23      ====        sub s9, a6, s7
                                                  30'd    6339    : data = 32'h    B60E4D93    ;    //    xori x27 x28 -1184      ====        xori s11, t3, -1184
                                                  30'd    6340    : data = 32'h    418C5013    ;    //    srai x0 x24 24      ====        srai zero, s8, 24
                                                  30'd    6341    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6342    : data = 32'h    3CC23493    ;    //    sltiu x9 x4 972      ====        sltiu s1, tp, 972
                                                  30'd    6343    : data = 32'h    8179B813    ;    //    sltiu x16 x19 -2025      ====        sltiu a6, s3, -2025
                                                  30'd    6344    : data = 32'h    15F30493    ;    //    addi x9 x6 351      ====        addi s1, t1, 351
                                                  30'd    6345    : data = 32'h    C47E8B13    ;    //    addi x22 x29 -953      ====        addi s6, t4, -953
                                                  30'd    6346    : data = 32'h    4057DB13    ;    //    srai x22 x15 5      ====        srai s6, a5, 5
                                                  30'd    6347    : data = 32'h    F3CA6293    ;    //    ori x5 x20 -196      ====        ori t0, s4, -196
                                                  30'd    6348    : data = 32'h    00A77AB3    ;    //    and x21 x14 x10      ====        and s5, a4, a0
                                                  30'd    6349    : data = 32'h    006E4FB3    ;    //    xor x31 x28 x6      ====        xor t6, t3, t1
                                                  30'd    6350    : data = 32'h    B46C3C13    ;    //    sltiu x24 x24 -1210      ====        sltiu s8, s8, -1210
                                                  30'd    6351    : data = 32'h    EEAC2A97    ;    //    auipc x21 977602      ====        auipc s5, 977602
                                                  30'd    6352    : data = 32'h    000202B3    ;    //    add x5 x4 x0      ====        add t0, tp, zero
                                                  30'd    6353    : data = 32'h    41B55713    ;    //    srai x14 x10 27      ====        srai a4, a0, 27
                                                  30'd    6354    : data = 32'h    01214BB3    ;    //    xor x23 x2 x18      ====        xor s7, sp, s2
                                                  30'd    6355    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6356    : data = 32'h    01AF26B3    ;    //    slt x13 x30 x26      ====        slt a3, t5, s10
                                                  30'd    6357    : data = 32'h    01997133    ;    //    and x2 x18 x25      ====        and sp, s2, s9
                                                  30'd    6358    : data = 32'h    D3208B13    ;    //    addi x22 x1 -718      ====        addi s6, ra, -718
                                                  30'd    6359    : data = 32'h    77BCC793    ;    //    xori x15 x25 1915      ====        xori a5, s9, 1915
                                                  30'd    6360    : data = 32'h    00703033    ;    //    sltu x0 x0 x7      ====        sltu zero, zero, t2
                                                  30'd    6361    : data = 32'h    01E4D913    ;    //    srli x18 x9 30      ====        srli s2, s1, 30
                                                  30'd    6362    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6363    : data = 32'h    01960DB3    ;    //    add x27 x12 x25      ====        add s11, a2, s9
                                                  30'd    6364    : data = 32'h    01308EB3    ;    //    add x29 x1 x19      ====        add t4, ra, s3
                                                  30'd    6365    : data = 32'h    F928F913    ;    //    andi x18 x17 -110      ====        andi s2, a7, -110
                                                  30'd    6366    : data = 32'h    0043D493    ;    //    srli x9 x7 4      ====        srli s1, t2, 4
                                                  30'd    6367    : data = 32'h    019E8833    ;    //    add x16 x29 x25      ====        add a6, t4, s9
                                                  30'd    6368    : data = 32'h    C14EA013    ;    //    slti x0 x29 -1004      ====        slti zero, t4, -1004
                                                  30'd    6369    : data = 32'h    4AD1E093    ;    //    ori x1 x3 1197      ====        ori ra, gp, 1197
                                                  30'd    6370    : data = 32'h    01E45633    ;    //    srl x12 x8 x30      ====        srl a2, s0, t5
                                                  30'd    6371    : data = 32'h    61472617    ;    //    auipc x12 398450      ====        auipc a2, 398450
                                                  30'd    6372    : data = 32'h    016148B3    ;    //    xor x17 x2 x22      ====        xor a7, sp, s6
                                                  30'd    6373    : data = 32'h    6CB0A037    ;    //    lui x0 445194      ====        lui zero, 445194
                                                  30'd    6374    : data = 32'h    014672B3    ;    //    and x5 x12 x20      ====        and t0, a2, s4
                                                  30'd    6375    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6376    : data = 32'h    0BE2AD93    ;    //    slti x27 x5 190      ====        slti s11, t0, 190
                                                  30'd    6377    : data = 32'h    00BBCD33    ;    //    xor x26 x23 x11      ====        xor s10, s7, a1
                                                  30'd    6378    : data = 32'h    00F682B3    ;    //    add x5 x13 x15      ====        add t0, a3, a5
                                                  30'd    6379    : data = 32'h    005E5293    ;    //    srli x5 x28 5      ====        srli t0, t3, 5
                                                  30'd    6380    : data = 32'h    0058BB33    ;    //    sltu x22 x17 x5      ====        sltu s6, a7, t0
                                                  30'd    6381    : data = 32'h    410987B3    ;    //    sub x15 x19 x16      ====        sub a5, s3, a6
                                                  30'd    6382    : data = 32'h    9B79E613    ;    //    ori x12 x19 -1609      ====        ori a2, s3, -1609
                                                  30'd    6383    : data = 32'h    41B3DA13    ;    //    srai x20 x7 27      ====        srai s4, t2, 27
                                                  30'd    6384    : data = 32'h    01551EB3    ;    //    sll x29 x10 x21      ====        sll t4, a0, s5
                                                  30'd    6385    : data = 32'h    01A2BA33    ;    //    sltu x20 x5 x26      ====        sltu s4, t0, s10
                                                  30'd    6386    : data = 32'h    00A52D33    ;    //    slt x26 x10 x10      ====        slt s10, a0, a0
                                                  30'd    6387    : data = 32'h    000261B3    ;    //    or x3 x4 x0      ====        or gp, tp, zero
                                                  30'd    6388    : data = 32'h    00DCDE13    ;    //    srli x28 x25 13      ====        srli t3, s9, 13
                                                  30'd    6389    : data = 32'h    1981C313    ;    //    xori x6 x3 408      ====        xori t1, gp, 408
                                                  30'd    6390    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6391    : data = 32'h    4029D713    ;    //    srai x14 x19 2      ====        srai a4, s3, 2
                                                  30'd    6392    : data = 32'h    09B6C093    ;    //    xori x1 x13 155      ====        xori ra, a3, 155
                                                  30'd    6393    : data = 32'h    00868433    ;    //    add x8 x13 x8      ====        add s0, a3, s0
                                                  30'd    6394    : data = 32'h    00025733    ;    //    srl x14 x4 x0      ====        srl a4, tp, zero
                                                  30'd    6395    : data = 32'h    00633D33    ;    //    sltu x26 x6 x6      ====        sltu s10, t1, t1
                                                  30'd    6396    : data = 32'h    40B48133    ;    //    sub x2 x9 x11      ====        sub sp, s1, a1
                                                  30'd    6397    : data = 32'h    B6C8C197    ;    //    auipc x3 748684      ====        auipc gp, 748684
                                                  30'd    6398    : data = 32'h    41185333    ;    //    sra x6 x16 x17      ====        sra t1, a6, a7
                                                  30'd    6399    : data = 32'h    00F28433    ;    //    add x8 x5 x15      ====        add s0, t0, a5
                                                  30'd    6400    : data = 32'h    41EA0433    ;    //    sub x8 x20 x30      ====        sub s0, s4, t5
                                                  30'd    6401    : data = 32'h    0B8ABB93    ;    //    sltiu x23 x21 184      ====        sltiu s7, s5, 184
                                                  30'd    6402    : data = 32'h    01FD5633    ;    //    srl x12 x26 x31      ====        srl a2, s10, t6
                                                  30'd    6403    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6404    : data = 32'h    00E31BB3    ;    //    sll x23 x6 x14      ====        sll s7, t1, a4
                                                  30'd    6405    : data = 32'h    2D9BE913    ;    //    ori x18 x23 729      ====        ori s2, s7, 729
                                                  30'd    6406    : data = 32'h    98C22F93    ;    //    slti x31 x4 -1652      ====        slti t6, tp, -1652
                                                  30'd    6407    : data = 32'h    00FB86B3    ;    //    add x13 x23 x15      ====        add a3, s7, a5
                                                  30'd    6408    : data = 32'h    405B5D13    ;    //    srai x26 x22 5      ====        srai s10, s6, 5
                                                  30'd    6409    : data = 32'h    C4E47013    ;    //    andi x0 x8 -946      ====        andi zero, s0, -946
                                                  30'd    6410    : data = 32'h    01E55C93    ;    //    srli x25 x10 30      ====        srli s9, a0, 30
                                                  30'd    6411    : data = 32'h    412DD813    ;    //    srai x16 x27 18      ====        srai a6, s11, 18
                                                  30'd    6412    : data = 32'h    D12BC013    ;    //    xori x0 x23 -750      ====        xori zero, s7, -750
                                                  30'd    6413    : data = 32'h    403B5E93    ;    //    srai x29 x22 3      ====        srai t4, s6, 3
                                                  30'd    6414    : data = 32'h    D1698E13    ;    //    addi x28 x19 -746      ====        addi t3, s3, -746
                                                  30'd    6415    : data = 32'h    82828097    ;    //    auipc x1 534568      ====        auipc ra, 534568
                                                  30'd    6416    : data = 32'h    29B7F313    ;    //    andi x6 x15 667      ====        andi t1, a5, 667
                                                  30'd    6417    : data = 32'h    0074B3B3    ;    //    sltu x7 x9 x7      ====        sltu t2, s1, t2
                                                  30'd    6418    : data = 32'h    1F19EC93    ;    //    ori x25 x19 497      ====        ori s9, s3, 497
                                                  30'd    6419    : data = 32'h    32E72297    ;    //    auipc x5 208498      ====        auipc t0, 208498
                                                  30'd    6420    : data = 32'h    00CFD093    ;    //    srli x1 x31 12      ====        srli ra, t6, 12
                                                  30'd    6421    : data = 32'h    E0D1CA93    ;    //    xori x21 x3 -499      ====        xori s5, gp, -499
                                                  30'd    6422    : data = 32'h    290E8493    ;    //    addi x9 x29 656      ====        addi s1, t4, 656
                                                  30'd    6423    : data = 32'h    00190C33    ;    //    add x24 x18 x1      ====        add s8, s2, ra
                                                  30'd    6424    : data = 32'h    00C51713    ;    //    slli x14 x10 12      ====        slli a4, a0, 12
                                                  30'd    6425    : data = 32'h    4FFC7093    ;    //    andi x1 x24 1279      ====        andi ra, s8, 1279
                                                  30'd    6426    : data = 32'h    2119BE13    ;    //    sltiu x28 x19 529      ====        sltiu t3, s3, 529
                                                  30'd    6427    : data = 32'h    018DA033    ;    //    slt x0 x27 x24      ====        slt zero, s11, s8
                                                  30'd    6428    : data = 32'h    00DF5E93    ;    //    srli x29 x30 13      ====        srli t4, t5, 13
                                                  30'd    6429    : data = 32'h    00D31093    ;    //    slli x1 x6 13      ====        slli ra, t1, 13
                                                  30'd    6430    : data = 32'h    0136CE33    ;    //    xor x28 x13 x19      ====        xor t3, a3, s3
                                                  30'd    6431    : data = 32'h    25F37813    ;    //    andi x16 x6 607      ====        andi a6, t1, 607
                                                  30'd    6432    : data = 32'h    35B43D13    ;    //    sltiu x26 x8 859      ====        sltiu s10, s0, 859
                                                  30'd    6433    : data = 32'h    00CA6833    ;    //    or x16 x20 x12      ====        or a6, s4, a2
                                                  30'd    6434    : data = 32'h    6F78F113    ;    //    andi x2 x17 1783      ====        andi sp, a7, 1783
                                                  30'd    6435    : data = 32'h    014D3933    ;    //    sltu x18 x26 x20      ====        sltu s2, s10, s4
                                                  30'd    6436    : data = 32'h    01925113    ;    //    srli x2 x4 25      ====        srli sp, tp, 25
                                                  30'd    6437    : data = 32'h    007A5EB3    ;    //    srl x29 x20 x7      ====        srl t4, s4, t2
                                                  30'd    6438    : data = 32'h    4544A837    ;    //    lui x16 283722      ====        lui a6, 283722
                                                  30'd    6439    : data = 32'h    4172DC93    ;    //    srai x25 x5 23      ====        srai s9, t0, 23
                                                  30'd    6440    : data = 32'h    0A3AE593    ;    //    ori x11 x21 163      ====        ori a1, s5, 163
                                                  30'd    6441    : data = 32'h    00BD1413    ;    //    slli x8 x26 11      ====        slli s0, s10, 11
                                                  30'd    6442    : data = 32'h    110B2693    ;    //    slti x13 x22 272      ====        slti a3, s6, 272
                                                  30'd    6443    : data = 32'h    40B586B3    ;    //    sub x13 x11 x11      ====        sub a3, a1, a1
                                                  30'd    6444    : data = 32'h    000AB0B3    ;    //    sltu x1 x21 x0      ====        sltu ra, s5, zero
                                                  30'd    6445    : data = 32'h    8F8520B7    ;    //    lui x1 587858      ====        lui ra, 587858
                                                  30'd    6446    : data = 32'h    01585833    ;    //    srl x16 x16 x21      ====        srl a6, a6, s5
                                                  30'd    6447    : data = 32'h    00099033    ;    //    sll x0 x19 x0      ====        sll zero, s3, zero
                                                  30'd    6448    : data = 32'h    00E82EB3    ;    //    slt x29 x16 x14      ====        slt t4, a6, a4
                                                  30'd    6449    : data = 32'h    01E3C1B3    ;    //    xor x3 x7 x30      ====        xor gp, t2, t5
                                                  30'd    6450    : data = 32'h    008DC633    ;    //    xor x12 x27 x8      ====        xor a2, s11, s0
                                                  30'd    6451    : data = 32'h    0019DD33    ;    //    srl x26 x19 x1      ====        srl s10, s3, ra
                                                  30'd    6452    : data = 32'h    75573D13    ;    //    sltiu x26 x14 1877      ====        sltiu s10, a4, 1877
                                                  30'd    6453    : data = 32'h    2FE7C193    ;    //    xori x3 x15 766      ====        xori gp, a5, 766
                                                  30'd    6454    : data = 32'h    1C0CE193    ;    //    ori x3 x25 448      ====        ori gp, s9, 448
                                                  30'd    6455    : data = 32'h    062FF637    ;    //    lui x12 25343      ====        lui a2, 25343
                                                  30'd    6456    : data = 32'h    4210EA13    ;    //    ori x20 x1 1057      ====        ori s4, ra, 1057
                                                  30'd    6457    : data = 32'h    9C550E93    ;    //    addi x29 x10 -1595      ====        addi t4, a0, -1595
                                                  30'd    6458    : data = 32'h    DAE78297    ;    //    auipc x5 896632      ====        auipc t0, 896632
                                                  30'd    6459    : data = 32'h    00F38CB3    ;    //    add x25 x7 x15      ====        add s9, t2, a5
                                                  30'd    6460    : data = 32'h    404CDD93    ;    //    srai x27 x25 4      ====        srai s11, s9, 4
                                                  30'd    6461    : data = 32'h    577EEC13    ;    //    ori x24 x29 1399      ====        ori s8, t4, 1399
                                                  30'd    6462    : data = 32'h    00D4D693    ;    //    srli x13 x9 13      ====        srli a3, s1, 13
                                                  30'd    6463    : data = 32'h    5531E713    ;    //    ori x14 x3 1363      ====        ori a4, gp, 1363
                                                  30'd    6464    : data = 32'h    AD083297    ;    //    auipc x5 708739      ====        auipc t0, 708739
                                                  30'd    6465    : data = 32'h    00381433    ;    //    sll x8 x16 x3      ====        sll s0, a6, gp
                                                  30'd    6466    : data = 32'h    00866633    ;    //    or x12 x12 x8      ====        or a2, a2, s0
                                                  30'd    6467    : data = 32'h    00795F93    ;    //    srli x31 x18 7      ====        srli t6, s2, 7
                                                  30'd    6468    : data = 32'h    4109D113    ;    //    srai x2 x19 16      ====        srai sp, s3, 16
                                                  30'd    6469    : data = 32'h    82170B13    ;    //    addi x22 x14 -2015      ====        addi s6, a4, -2015
                                                  30'd    6470    : data = 32'h    5EA0C993    ;    //    xori x19 x1 1514      ====        xori s3, ra, 1514
                                                  30'd    6471    : data = 32'h    00583833    ;    //    sltu x16 x16 x5      ====        sltu a6, a6, t0
                                                  30'd    6472    : data = 32'h    40DB5393    ;    //    srai x7 x22 13      ====        srai t2, s6, 13
                                                  30'd    6473    : data = 32'h    4422B193    ;    //    sltiu x3 x5 1090      ====        sltiu gp, t0, 1090
                                                  30'd    6474    : data = 32'h    1AF13593    ;    //    sltiu x11 x2 431      ====        sltiu a1, sp, 431
                                                  30'd    6475    : data = 32'h    41B6D913    ;    //    srai x18 x13 27      ====        srai s2, a3, 27
                                                  30'd    6476    : data = 32'h    014BD633    ;    //    srl x12 x23 x20      ====        srl a2, s7, s4
                                                  30'd    6477    : data = 32'h    E6F2F813    ;    //    andi x16 x5 -401      ====        andi a6, t0, -401
                                                  30'd    6478    : data = 32'h    0059D713    ;    //    srli x14 x19 5      ====        srli a4, s3, 5
                                                  30'd    6479    : data = 32'h    018FB833    ;    //    sltu x16 x31 x24      ====        sltu a6, t6, s8
                                                  30'd    6480    : data = 32'h    01E228B3    ;    //    slt x17 x4 x30      ====        slt a7, tp, t5
                                                  30'd    6481    : data = 32'h    00C97BB3    ;    //    and x23 x18 x12      ====        and s7, s2, a2
                                                  30'd    6482    : data = 32'h    40815393    ;    //    srai x7 x2 8      ====        srai t2, sp, 8
                                                  30'd    6483    : data = 32'h    FD052C13    ;    //    slti x24 x10 -48      ====        slti s8, a0, -48
                                                  30'd    6484    : data = 32'h    01228E33    ;    //    add x28 x5 x18      ====        add t3, t0, s2
                                                  30'd    6485    : data = 32'h    0C18FC13    ;    //    andi x24 x17 193      ====        andi s8, a7, 193
                                                  30'd    6486    : data = 32'h    012F1093    ;    //    slli x1 x30 18      ====        slli ra, t5, 18
                                                  30'd    6487    : data = 32'h    D2AF89B7    ;    //    lui x19 862968      ====        lui s3, 862968
                                                  30'd    6488    : data = 32'h    41C05693    ;    //    srai x13 x0 28      ====        srai a3, zero, 28
                                                  30'd    6489    : data = 32'h    97EA2813    ;    //    slti x16 x20 -1666      ====        slti a6, s4, -1666
                                                  30'd    6490    : data = 32'h    01417C33    ;    //    and x24 x2 x20      ====        and s8, sp, s4
                                                  30'd    6491    : data = 32'h    005D4C33    ;    //    xor x24 x26 x5      ====        xor s8, s10, t0
                                                  30'd    6492    : data = 32'h    409ED133    ;    //    sra x2 x29 x9      ====        sra sp, t4, s1
                                                  30'd    6493    : data = 32'h    001CFB33    ;    //    and x22 x25 x1      ====        and s6, s9, ra
                                                  30'd    6494    : data = 32'h    8E2AA313    ;    //    slti x6 x21 -1822      ====        slti t1, s5, -1822
                                                  30'd    6495    : data = 32'h    401FDA33    ;    //    sra x20 x31 x1      ====        sra s4, t6, ra
                                                  30'd    6496    : data = 32'h    0006A733    ;    //    slt x14 x13 x0      ====        slt a4, a3, zero
                                                  30'd    6497    : data = 32'h    01D35093    ;    //    srli x1 x6 29      ====        srli ra, t1, 29
                                                  30'd    6498    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6499    : data = 32'h    00E81A13    ;    //    slli x20 x16 14      ====        slli s4, a6, 14
                                                  30'd    6500    : data = 32'h    00BF1E13    ;    //    slli x28 x30 11      ====        slli t3, t5, 11
                                                  30'd    6501    : data = 32'h    41890033    ;    //    sub x0 x18 x24      ====        sub zero, s2, s8
                                                  30'd    6502    : data = 32'h    013586B3    ;    //    add x13 x11 x19      ====        add a3, a1, s3
                                                  30'd    6503    : data = 32'h    41798433    ;    //    sub x8 x19 x23      ====        sub s0, s3, s7
                                                  30'd    6504    : data = 32'h    00F86DB3    ;    //    or x27 x16 x15      ====        or s11, a6, a5
                                                  30'd    6505    : data = 32'h    00B41833    ;    //    sll x16 x8 x11      ====        sll a6, s0, a1
                                                  30'd    6506    : data = 32'h    0137B433    ;    //    sltu x8 x15 x19      ====        sltu s0, a5, s3
                                                  30'd    6507    : data = 32'h    00309633    ;    //    sll x12 x1 x3      ====        sll a2, ra, gp
                                                  30'd    6508    : data = 32'h    9C34B113    ;    //    sltiu x2 x9 -1597      ====        sltiu sp, s1, -1597
                                                  30'd    6509    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6510    : data = 32'h    40E387B3    ;    //    sub x15 x7 x14      ====        sub a5, t2, a4
                                                  30'd    6511    : data = 32'h    014BCDB3    ;    //    xor x27 x23 x20      ====        xor s11, s7, s4
                                                  30'd    6512    : data = 32'h    000407B3    ;    //    add x15 x8 x0      ====        add a5, s0, zero
                                                  30'd    6513    : data = 32'h    01A03CB3    ;    //    sltu x25 x0 x26      ====        sltu s9, zero, s10
                                                  30'd    6514    : data = 32'h    001CC933    ;    //    xor x18 x25 x1      ====        xor s2, s9, ra
                                                  30'd    6515    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6516    : data = 32'h    0EF8AF93    ;    //    slti x31 x17 239      ====        slti t6, a7, 239
                                                  30'd    6517    : data = 32'h    004F5E33    ;    //    srl x28 x30 x4      ====        srl t3, t5, tp
                                                  30'd    6518    : data = 32'h    00CCC5B3    ;    //    xor x11 x25 x12      ====        xor a1, s9, a2
                                                  30'd    6519    : data = 32'h    00171093    ;    //    slli x1 x14 1      ====        slli ra, a4, 1
                                                  30'd    6520    : data = 32'h    381BCC13    ;    //    xori x24 x23 897      ====        xori s8, s7, 897
                                                  30'd    6521    : data = 32'h    C17D3E13    ;    //    sltiu x28 x26 -1001      ====        sltiu t3, s10, -1001
                                                  30'd    6522    : data = 32'h    6B293D13    ;    //    sltiu x26 x18 1714      ====        sltiu s10, s2, 1714
                                                  30'd    6523    : data = 32'h    41D55733    ;    //    sra x14 x10 x29      ====        sra a4, a0, t4
                                                  30'd    6524    : data = 32'h    27286413    ;    //    ori x8 x16 626      ====        ori s0, a6, 626
                                                  30'd    6525    : data = 32'h    403B5E13    ;    //    srai x28 x22 3      ====        srai t3, s6, 3
                                                  30'd    6526    : data = 32'h    416FD433    ;    //    sra x8 x31 x22      ====        sra s0, t6, s6
                                                  30'd    6527    : data = 32'h    23E33093    ;    //    sltiu x1 x6 574      ====        sltiu ra, t1, 574
                                                  30'd    6528    : data = 32'h    2462E193    ;    //    ori x3 x5 582      ====        ori gp, t0, 582
                                                  30'd    6529    : data = 32'h    00140733    ;    //    add x14 x8 x1      ====        add a4, s0, ra
                                                  30'd    6530    : data = 32'h    0092DA33    ;    //    srl x20 x5 x9      ====        srl s4, t0, s1
                                                  30'd    6531    : data = 32'h    49CDE913    ;    //    ori x18 x27 1180      ====        ori s2, s11, 1180
                                                  30'd    6532    : data = 32'h    014A76B3    ;    //    and x13 x20 x20      ====        and a3, s4, s4
                                                  30'd    6533    : data = 32'h    1C24EA17    ;    //    auipc x20 115278      ====        auipc s4, 115278
                                                  30'd    6534    : data = 32'h    86DAA493    ;    //    slti x9 x21 -1939      ====        slti s1, s5, -1939
                                                  30'd    6535    : data = 32'h    00ECF5B3    ;    //    and x11 x25 x14      ====        and a1, s9, a4
                                                  30'd    6536    : data = 32'h    00CAB2B3    ;    //    sltu x5 x21 x12      ====        sltu t0, s5, a2
                                                  30'd    6537    : data = 32'h    00B69093    ;    //    slli x1 x13 11      ====        slli ra, a3, 11
                                                  30'd    6538    : data = 32'h    41D45C33    ;    //    sra x24 x8 x29      ====        sra s8, s0, t4
                                                  30'd    6539    : data = 32'h    F407A193    ;    //    slti x3 x15 -192      ====        slti gp, a5, -192
                                                  30'd    6540    : data = 32'h    01B3D633    ;    //    srl x12 x7 x27      ====        srl a2, t2, s11
                                                  30'd    6541    : data = 32'h    00E69613    ;    //    slli x12 x13 14      ====        slli a2, a3, 14
                                                  30'd    6542    : data = 32'h    017DE433    ;    //    or x8 x27 x23      ====        or s0, s11, s7
                                                  30'd    6543    : data = 32'h    011DCCB3    ;    //    xor x25 x27 x17      ====        xor s9, s11, a7
                                                  30'd    6544    : data = 32'h    0191D013    ;    //    srli x0 x3 25      ====        srli zero, gp, 25
                                                  30'd    6545    : data = 32'h    01C39E93    ;    //    slli x29 x7 28      ====        slli t4, t2, 28
                                                  30'd    6546    : data = 32'h    DF5A5B97    ;    //    auipc x23 914853      ====        auipc s7, 914853
                                                  30'd    6547    : data = 32'h    406AD013    ;    //    srai x0 x21 6      ====        srai zero, s5, 6
                                                  30'd    6548    : data = 32'h    4129D033    ;    //    sra x0 x19 x18      ====        sra zero, s3, s2
                                                  30'd    6549    : data = 32'h    69563E13    ;    //    sltiu x28 x12 1685      ====        sltiu t3, a2, 1685
                                                  30'd    6550    : data = 32'h    01F8B733    ;    //    sltu x14 x17 x31      ====        sltu a4, a7, t6
                                                  30'd    6551    : data = 32'h    0029BD33    ;    //    sltu x26 x19 x2      ====        sltu s10, s3, sp
                                                  30'd    6552    : data = 32'h    F0020A13    ;    //    addi x20 x4 -256      ====        addi s4, tp, -256
                                                  30'd    6553    : data = 32'h    01F8F7B3    ;    //    and x15 x17 x31      ====        and a5, a7, t6
                                                  30'd    6554    : data = 32'h    0F9AAE93    ;    //    slti x29 x21 249      ====        slti t4, s5, 249
                                                  30'd    6555    : data = 32'h    0030CBB3    ;    //    xor x23 x1 x3      ====        xor s7, ra, gp
                                                  30'd    6556    : data = 32'h    00FBB7B3    ;    //    sltu x15 x23 x15      ====        sltu a5, s7, a5
                                                  30'd    6557    : data = 32'h    01D3EB33    ;    //    or x22 x7 x29      ====        or s6, t2, t4
                                                  30'd    6558    : data = 32'h    412350B3    ;    //    sra x1 x6 x18      ====        sra ra, t1, s2
                                                  30'd    6559    : data = 32'h    B0B88D13    ;    //    addi x26 x17 -1269      ====        addi s10, a7, -1269
                                                  30'd    6560    : data = 32'h    019B5BB3    ;    //    srl x23 x22 x25      ====        srl s7, s6, s9
                                                  30'd    6561    : data = 32'h    8EAD6397    ;    //    auipc x7 584406      ====        auipc t2, 584406
                                                  30'd    6562    : data = 32'h    DB8FBE13    ;    //    sltiu x28 x31 -584      ====        sltiu t3, t6, -584
                                                  30'd    6563    : data = 32'h    F73B5497    ;    //    auipc x9 1012661      ====        auipc s1, 1012661
                                                  30'd    6564    : data = 32'h    249366B7    ;    //    lui x13 149814      ====        lui a3, 149814
                                                  30'd    6565    : data = 32'h    01F0B0B3    ;    //    sltu x1 x1 x31      ====        sltu ra, ra, t6
                                                  30'd    6566    : data = 32'h    019B35B3    ;    //    sltu x11 x22 x25      ====        sltu a1, s6, s9
                                                  30'd    6567    : data = 32'h    00F758B3    ;    //    srl x17 x14 x15      ====        srl a7, a4, a5
                                                  30'd    6568    : data = 32'h    D5496D13    ;    //    ori x26 x18 -684      ====        ori s10, s2, -684
                                                  30'd    6569    : data = 32'h    01F20633    ;    //    add x12 x4 x31      ====        add a2, tp, t6
                                                  30'd    6570    : data = 32'h    7B3F0993    ;    //    addi x19 x30 1971      ====        addi s3, t5, 1971
                                                  30'd    6571    : data = 32'h    00EA4B33    ;    //    xor x22 x20 x14      ====        xor s6, s4, a4
                                                  30'd    6572    : data = 32'h    00C0D993    ;    //    srli x19 x1 12      ====        srli s3, ra, 12
                                                  30'd    6573    : data = 32'h    40F75093    ;    //    srai x1 x14 15      ====        srai ra, a4, 15
                                                  30'd    6574    : data = 32'h    00BAA433    ;    //    slt x8 x21 x11      ====        slt s0, s5, a1
                                                  30'd    6575    : data = 32'h    00524FB3    ;    //    xor x31 x4 x5      ====        xor t6, tp, t0
                                                  30'd    6576    : data = 32'h    E2E6C417    ;    //    auipc x8 929388      ====        auipc s0, 929388
                                                  30'd    6577    : data = 32'h    01836133    ;    //    or x2 x6 x24      ====        or sp, t1, s8
                                                  30'd    6578    : data = 32'h    044FB813    ;    //    sltiu x16 x31 68      ====        sltiu a6, t6, 68
                                                  30'd    6579    : data = 32'h    00D4DD33    ;    //    srl x26 x9 x13      ====        srl s10, s1, a3
                                                  30'd    6580    : data = 32'h    014D1313    ;    //    slli x6 x26 20      ====        slli t1, s10, 20
                                                  30'd    6581    : data = 32'h    409B4C93    ;    //    xori x25 x22 1033      ====        xori s9, s6, 1033
                                                  30'd    6582    : data = 32'h    8E278B93    ;    //    addi x23 x15 -1822      ====        addi s7, a5, -1822
                                                  30'd    6583    : data = 32'h    1AB14313    ;    //    xori x6 x2 427      ====        xori t1, sp, 427
                                                  30'd    6584    : data = 32'h    09E05437    ;    //    lui x8 40453      ====        lui s0, 40453
                                                  30'd    6585    : data = 32'h    406E88B3    ;    //    sub x17 x29 x6      ====        sub a7, t4, t1
                                                  30'd    6586    : data = 32'h    5DAE8BB7    ;    //    lui x23 383720      ====        lui s7, 383720
                                                  30'd    6587    : data = 32'h    9A6FA113    ;    //    slti x2 x31 -1626      ====        slti sp, t6, -1626
                                                  30'd    6588    : data = 32'h    012A6DB3    ;    //    or x27 x20 x18      ====        or s11, s4, s2
                                                  30'd    6589    : data = 32'h    017B20B3    ;    //    slt x1 x22 x23      ====        slt ra, s6, s7
                                                  30'd    6590    : data = 32'h    417104B3    ;    //    sub x9 x2 x23      ====        sub s1, sp, s7
                                                  30'd    6591    : data = 32'h    BA97B993    ;    //    sltiu x19 x15 -1111      ====        sltiu s3, a5, -1111
                                                  30'd    6592    : data = 32'h    A8419117    ;    //    auipc x2 689177      ====        auipc sp, 689177
                                                  30'd    6593    : data = 32'h    00B7F7B3    ;    //    and x15 x15 x11      ====        and a5, a5, a1
                                                  30'd    6594    : data = 32'h    96DECC93    ;    //    xori x25 x29 -1683      ====        xori s9, t4, -1683
                                                  30'd    6595    : data = 32'h    F245CBB7    ;    //    lui x23 992348      ====        lui s7, 992348
                                                  30'd    6596    : data = 32'h    000BE0B3    ;    //    or x1 x23 x0      ====        or ra, s7, zero
                                                  30'd    6597    : data = 32'h    00027B33    ;    //    and x22 x4 x0      ====        and s6, tp, zero
                                                  30'd    6598    : data = 32'h    41945C33    ;    //    sra x24 x8 x25      ====        sra s8, s0, s9
                                                  30'd    6599    : data = 32'h    00DE73B3    ;    //    and x7 x28 x13      ====        and t2, t3, a3
                                                  30'd    6600    : data = 32'h    00C7A733    ;    //    slt x14 x15 x12      ====        slt a4, a5, a2
                                                  30'd    6601    : data = 32'h    00D2C133    ;    //    xor x2 x5 x13      ====        xor sp, t0, a3
                                                  30'd    6602    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6603    : data = 32'h    DB543017    ;    //    auipc x0 898371      ====        auipc zero, 898371
                                                  30'd    6604    : data = 32'h    7DE7BD93    ;    //    sltiu x27 x15 2014      ====        sltiu s11, a5, 2014
                                                  30'd    6605    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6606    : data = 32'h    68EB3D13    ;    //    sltiu x26 x22 1678      ====        sltiu s10, s6, 1678
                                                  30'd    6607    : data = 32'h    42392713    ;    //    slti x14 x18 1059      ====        slti a4, s2, 1059
                                                  30'd    6608    : data = 32'h    B33A6C93    ;    //    ori x25 x20 -1229      ====        ori s9, s4, -1229
                                                  30'd    6609    : data = 32'h    018AB5B3    ;    //    sltu x11 x21 x24      ====        sltu a1, s5, s8
                                                  30'd    6610    : data = 32'h    00CD93B3    ;    //    sll x7 x27 x12      ====        sll t2, s11, a2
                                                  30'd    6611    : data = 32'h    01851813    ;    //    slli x16 x10 24      ====        slli a6, a0, 24
                                                  30'd    6612    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6613    : data = 32'h    16386893    ;    //    ori x17 x16 355      ====        ori a7, a6, 355
                                                  30'd    6614    : data = 32'h    00006633    ;    //    or x12 x0 x0      ====        or a2, zero, zero
                                                  30'd    6615    : data = 32'h    00011E33    ;    //    sll x28 x2 x0      ====        sll t3, sp, zero
                                                  30'd    6616    : data = 32'h    40580033    ;    //    sub x0 x16 x5      ====        sub zero, a6, t0
                                                  30'd    6617    : data = 32'h    00000113    ;    //    addi x2 x0 0      ====        li sp, 0x0 #start riscv_int_numeric_corner_stream_38
                                                  30'd    6618    : data = 32'h    800000B7    ;    //    lui x1 524288      ====        li ra, 0x80000000
                                                  30'd    6619    : data = 32'h    00008093    ;    //    addi x1 x1 0      ====        li ra, 0x80000000
                                                  30'd    6620    : data = 32'h    85AA8AB7    ;    //    lui x21 547496      ====        li s5, 0x85aa82b1
                                                  30'd    6621    : data = 32'h    2B1A8A93    ;    //    addi x21 x21 689      ====        li s5, 0x85aa82b1
                                                  30'd    6622    : data = 32'h    00000C13    ;    //    addi x24 x0 0      ====        li s8, 0x0
                                                  30'd    6623    : data = 32'h    748E8FB7    ;    //    lui x31 477416      ====        li t6, 0x748e7ccb
                                                  30'd    6624    : data = 32'h    CCBF8F93    ;    //    addi x31 x31 -821      ====        li t6, 0x748e7ccb
                                                  30'd    6625    : data = 32'h    800004B7    ;    //    lui x9 524288      ====        li s1, 0x80000000
                                                  30'd    6626    : data = 32'h    00048493    ;    //    addi x9 x9 0      ====        li s1, 0x80000000
                                                  30'd    6627    : data = 32'h    017EDB37    ;    //    lui x22 6125      ====        li s6, 0x17ed7a0
                                                  30'd    6628    : data = 32'h    7A0B0B13    ;    //    addi x22 x22 1952      ====        li s6, 0x17ed7a0
                                                  30'd    6629    : data = 32'h    FFF00D93    ;    //    addi x27 x0 -1      ====        li s11, 0xffffffff
                                                  30'd    6630    : data = 32'h    74F27BB7    ;    //    lui x23 479015      ====        li s7, 0x74f27535
                                                  30'd    6631    : data = 32'h    535B8B93    ;    //    addi x23 x23 1333      ====        li s7, 0x74f27535
                                                  30'd    6632    : data = 32'h    FFF00193    ;    //    addi x3 x0 -1      ====        li gp, 0xffffffff
                                                  30'd    6633    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6634    : data = 32'h    402A84B3    ;    //    sub x9 x21 x2      ====        sub s1, s5, sp
                                                  30'd    6635    : data = 32'h    C36EB1B7    ;    //    lui x3 800491      ====        lui gp, 800491
                                                  30'd    6636    : data = 32'h    837C0A93    ;    //    addi x21 x24 -1993      ====        addi s5, s8, -1993
                                                  30'd    6637    : data = 32'h    C58A4C17    ;    //    auipc x24 809124      ====        auipc s8, 809124
                                                  30'd    6638    : data = 32'h    4AD6E117    ;    //    auipc x2 306542      ====        auipc sp, 306542
                                                  30'd    6639    : data = 32'h    402B0BB3    ;    //    sub x23 x22 x2      ====        sub s7, s6, sp
                                                  30'd    6640    : data = 32'h    009184B3    ;    //    add x9 x3 x9      ====        add s1, gp, s1
                                                  30'd    6641    : data = 32'h    E1E08113    ;    //    addi x2 x1 -482      ====        addi sp, ra, -482
                                                  30'd    6642    : data = 32'h    416F8B33    ;    //    sub x22 x31 x22      ====        sub s6, t6, s6
                                                  30'd    6643    : data = 32'h    26630B97    ;    //    auipc x23 157232      ====        auipc s7, 157232
                                                  30'd    6644    : data = 32'h    C6D59117    ;    //    auipc x2 814425      ====        auipc sp, 814425
                                                  30'd    6645    : data = 32'h    FC64DA97    ;    //    auipc x21 1033805      ====        auipc s5, 1033805
                                                  30'd    6646    : data = 32'h    6B7D8493    ;    //    addi x9 x27 1719      ====        addi s1, s11, 1719
                                                  30'd    6647    : data = 32'h    5AD18B17    ;    //    auipc x22 371992      ====        auipc s6, 371992
                                                  30'd    6648    : data = 32'h    709040EF    ;    //    jal x1 20232      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_38
                                                  30'd    6649    : data = 32'h    FB8A8993    ;    //    addi x19 x21 -72      ====        addi s3, s5, -72
                                                  30'd    6650    : data = 32'h    A7780013    ;    //    addi x0 x16 -1417      ====        addi zero, a6, -1417
                                                  30'd    6651    : data = 32'h    5837E193    ;    //    ori x3 x15 1411      ====        ori gp, a5, 1411
                                                  30'd    6652    : data = 32'h    0055B333    ;    //    sltu x6 x11 x5      ====        sltu t1, a1, t0
                                                  30'd    6653    : data = 32'h    413887B3    ;    //    sub x15 x17 x19      ====        sub a5, a7, s3
                                                  30'd    6654    : data = 32'h    C0AD8C13    ;    //    addi x24 x27 -1014      ====        addi s8, s11, -1014
                                                  30'd    6655    : data = 32'h    00039913    ;    //    slli x18 x7 0      ====        slli s2, t2, 0
                                                  30'd    6656    : data = 32'h    8A05E413    ;    //    ori x8 x11 -1888      ====        ori s0, a1, -1888
                                                  30'd    6657    : data = 32'h    01A53133    ;    //    sltu x2 x10 x26      ====        sltu sp, a0, s10
                                                  30'd    6658    : data = 32'h    403D80B3    ;    //    sub x1 x27 x3      ====        sub ra, s11, gp
                                                  30'd    6659    : data = 32'h    757A8313    ;    //    addi x6 x21 1879      ====        addi t1, s5, 1879
                                                  30'd    6660    : data = 32'h    F5A3A1B7    ;    //    lui x3 1006138      ====        lui gp, 1006138
                                                  30'd    6661    : data = 32'h    466F0293    ;    //    addi x5 x30 1126      ====        addi t0, t5, 1126
                                                  30'd    6662    : data = 32'h    9C5682B7    ;    //    lui x5 640360      ====        lui t0, 640360
                                                  30'd    6663    : data = 32'h    4449E713    ;    //    ori x14 x19 1092      ====        ori a4, s3, 1092
                                                  30'd    6664    : data = 32'h    01F407B3    ;    //    add x15 x8 x31      ====        add a5, s0, t6
                                                  30'd    6665    : data = 32'h    4D103893    ;    //    sltiu x17 x0 1233      ====        sltiu a7, zero, 1233
                                                  30'd    6666    : data = 32'h    BFEBB097    ;    //    auipc x1 786107      ====        auipc ra, 786107
                                                  30'd    6667    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6668    : data = 32'h    00E7EAB3    ;    //    or x21 x15 x14      ====        or s5, a5, a4
                                                  30'd    6669    : data = 32'h    11ABAC93    ;    //    slti x25 x23 282      ====        slti s9, s7, 282
                                                  30'd    6670    : data = 32'h    013D5193    ;    //    srli x3 x26 19      ====        srli gp, s10, 19
                                                  30'd    6671    : data = 32'h    00E2EAB3    ;    //    or x21 x5 x14      ====        or s5, t0, a4
                                                  30'd    6672    : data = 32'h    01425D13    ;    //    srli x26 x4 20      ====        srli s10, tp, 20
                                                  30'd    6673    : data = 32'h    0B1E6E13    ;    //    ori x28 x28 177      ====        ori t3, t3, 177
                                                  30'd    6674    : data = 32'h    00DABC33    ;    //    sltu x24 x21 x13      ====        sltu s8, s5, a3
                                                  30'd    6675    : data = 32'h    000B03B3    ;    //    add x7 x22 x0      ====        add t2, s6, zero
                                                  30'd    6676    : data = 32'h    99FB9C17    ;    //    auipc x24 630713      ====        auipc s8, 630713
                                                  30'd    6677    : data = 32'h    416683B3    ;    //    sub x7 x13 x22      ====        sub t2, a3, s6
                                                  30'd    6678    : data = 32'h    00055593    ;    //    srli x11 x10 0      ====        srli a1, a0, 0
                                                  30'd    6679    : data = 32'h    00F238B3    ;    //    sltu x17 x4 x15      ====        sltu a7, tp, a5
                                                  30'd    6680    : data = 32'h    7E108C13    ;    //    addi x24 x1 2017      ====        addi s8, ra, 2017
                                                  30'd    6681    : data = 32'h    01F68433    ;    //    add x8 x13 x31      ====        add s0, a3, t6
                                                  30'd    6682    : data = 32'h    0067E7B3    ;    //    or x15 x15 x6      ====        or a5, a5, t1
                                                  30'd    6683    : data = 32'h    01F7D5B3    ;    //    srl x11 x15 x31      ====        srl a1, a5, t6
                                                  30'd    6684    : data = 32'h    41ECDBB3    ;    //    sra x23 x25 x30      ====        sra s7, s9, t5
                                                  30'd    6685    : data = 32'h    00195013    ;    //    srli x0 x18 1      ====        srli zero, s2, 1
                                                  30'd    6686    : data = 32'h    01809C93    ;    //    slli x25 x1 24      ====        slli s9, ra, 24
                                                  30'd    6687    : data = 32'h    01C52733    ;    //    slt x14 x10 x28      ====        slt a4, a0, t3
                                                  30'd    6688    : data = 32'h    1F5D8493    ;    //    addi x9 x27 501      ====        addi s1, s11, 501
                                                  30'd    6689    : data = 32'h    00555B13    ;    //    srli x22 x10 5      ====        srli s6, a0, 5
                                                  30'd    6690    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6691    : data = 32'h    01385D93    ;    //    srli x27 x16 19      ====        srli s11, a6, 19
                                                  30'd    6692    : data = 32'h    703D3717    ;    //    auipc x14 459731      ====        auipc a4, 459731
                                                  30'd    6693    : data = 32'h    01856EB3    ;    //    or x29 x10 x24      ====        or t4, a0, s8
                                                  30'd    6694    : data = 32'h    00FA37B3    ;    //    sltu x15 x20 x15      ====        sltu a5, s4, a5
                                                  30'd    6695    : data = 32'h    7C78F593    ;    //    andi x11 x17 1991      ====        andi a1, a7, 1991
                                                  30'd    6696    : data = 32'h    40175113    ;    //    srai x2 x14 1      ====        srai sp, a4, 1
                                                  30'd    6697    : data = 32'h    002701B3    ;    //    add x3 x14 x2      ====        add gp, a4, sp
                                                  30'd    6698    : data = 32'h    2F63B793    ;    //    sltiu x15 x7 758      ====        sltiu a5, t2, 758
                                                  30'd    6699    : data = 32'h    40655A33    ;    //    sra x20 x10 x6      ====        sra s4, a0, t1
                                                  30'd    6700    : data = 32'h    A0DA2337    ;    //    lui x6 658850      ====        lui t1, 658850
                                                  30'd    6701    : data = 32'h    081C6837    ;    //    lui x16 33222      ====        lui a6, 33222
                                                  30'd    6702    : data = 32'h    01C3F433    ;    //    and x8 x7 x28      ====        and s0, t2, t3
                                                  30'd    6703    : data = 32'h    E7D70B13    ;    //    addi x22 x14 -387      ====        addi s6, a4, -387
                                                  30'd    6704    : data = 32'h    0135F633    ;    //    and x12 x11 x19      ====        and a2, a1, s3
                                                  30'd    6705    : data = 32'h    7AB7F713    ;    //    andi x14 x15 1963      ====        andi a4, a5, 1963
                                                  30'd    6706    : data = 32'h    00501DB3    ;    //    sll x27 x0 x5      ====        sll s11, zero, t0
                                                  30'd    6707    : data = 32'h    00BBDB13    ;    //    srli x22 x23 11      ====        srli s6, s7, 11
                                                  30'd    6708    : data = 32'h    01531413    ;    //    slli x8 x6 21      ====        slli s0, t1, 21
                                                  30'd    6709    : data = 32'h    012DDA93    ;    //    srli x21 x27 18      ====        srli s5, s11, 18
                                                  30'd    6710    : data = 32'h    86714393    ;    //    xori x7 x2 -1945      ====        xori t2, sp, -1945
                                                  30'd    6711    : data = 32'h    015117B3    ;    //    sll x15 x2 x21      ====        sll a5, sp, s5
                                                  30'd    6712    : data = 32'h    006529B3    ;    //    slt x19 x10 x6      ====        slt s3, a0, t1
                                                  30'd    6713    : data = 32'h    01375CB3    ;    //    srl x25 x14 x19      ====        srl s9, a4, s3
                                                  30'd    6714    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6715    : data = 32'h    C6783713    ;    //    sltiu x14 x16 -921      ====        sltiu a4, a6, -921
                                                  30'd    6716    : data = 32'h    007C6633    ;    //    or x12 x24 x7      ====        or a2, s8, t2
                                                  30'd    6717    : data = 32'h    018D5A33    ;    //    srl x20 x26 x24      ====        srl s4, s10, s8
                                                  30'd    6718    : data = 32'h    F1570393    ;    //    addi x7 x14 -235      ====        addi t2, a4, -235
                                                  30'd    6719    : data = 32'h    01CCB833    ;    //    sltu x16 x25 x28      ====        sltu a6, s9, t3
                                                  30'd    6720    : data = 32'h    01702B33    ;    //    slt x22 x0 x23      ====        slt s6, zero, s7
                                                  30'd    6721    : data = 32'h    434F15B7    ;    //    lui x11 275697      ====        lui a1, 275697
                                                  30'd    6722    : data = 32'h    B046A293    ;    //    slti x5 x13 -1276      ====        slti t0, a3, -1276
                                                  30'd    6723    : data = 32'h    41C78FB3    ;    //    sub x31 x15 x28      ====        sub t6, a5, t3
                                                  30'd    6724    : data = 32'h    4031D6B3    ;    //    sra x13 x3 x3      ====        sra a3, gp, gp
                                                  30'd    6725    : data = 32'h    01215E13    ;    //    srli x28 x2 18      ====        srli t3, sp, 18
                                                  30'd    6726    : data = 32'h    40DE02B3    ;    //    sub x5 x28 x13      ====        sub t0, t3, a3
                                                  30'd    6727    : data = 32'h    6186A113    ;    //    slti x2 x13 1560      ====        slti sp, a3, 1560
                                                  30'd    6728    : data = 32'h    017C16B3    ;    //    sll x13 x24 x23      ====        sll a3, s8, s7
                                                  30'd    6729    : data = 32'h    448E0B93    ;    //    addi x23 x28 1096      ====        addi s7, t3, 1096
                                                  30'd    6730    : data = 32'h    B6F6AE13    ;    //    slti x28 x13 -1169      ====        slti t3, a3, -1169
                                                  30'd    6731    : data = 32'h    000AC733    ;    //    xor x14 x21 x0      ====        xor a4, s5, zero
                                                  30'd    6732    : data = 32'h    7FAEA793    ;    //    slti x15 x29 2042      ====        slti a5, t4, 2042
                                                  30'd    6733    : data = 32'h    41965693    ;    //    srai x13 x12 25      ====        srai a3, a2, 25
                                                  30'd    6734    : data = 32'h    00753D33    ;    //    sltu x26 x10 x7      ====        sltu s10, a0, t2
                                                  30'd    6735    : data = 32'h    25890E37    ;    //    lui x28 153744      ====        lui t3, 153744
                                                  30'd    6736    : data = 32'h    01BA6B33    ;    //    or x22 x20 x27      ====        or s6, s4, s11
                                                  30'd    6737    : data = 32'h    01F8DD93    ;    //    srli x27 x17 31      ====        srli s11, a7, 31
                                                  30'd    6738    : data = 32'h    41A182B3    ;    //    sub x5 x3 x26      ====        sub t0, gp, s10
                                                  30'd    6739    : data = 32'h    0003D3B3    ;    //    srl x7 x7 x0      ====        srl t2, t2, zero
                                                  30'd    6740    : data = 32'h    ED900113    ;    //    addi x2 x0 -295      ====        addi sp, zero, -295
                                                  30'd    6741    : data = 32'h    405403B3    ;    //    sub x7 x8 x5      ====        sub t2, s0, t0
                                                  30'd    6742    : data = 32'h    0064E6B3    ;    //    or x13 x9 x6      ====        or a3, s1, t1
                                                  30'd    6743    : data = 32'h    00BCAFB3    ;    //    slt x31 x25 x11      ====        slt t6, s9, a1
                                                  30'd    6744    : data = 32'h    110FE037    ;    //    lui x0 69886      ====        lui zero, 69886
                                                  30'd    6745    : data = 32'h    010DCD33    ;    //    xor x26 x27 x16      ====        xor s10, s11, a6
                                                  30'd    6746    : data = 32'h    41C5D3B3    ;    //    sra x7 x11 x28      ====        sra t2, a1, t3
                                                  30'd    6747    : data = 32'h    403FDF93    ;    //    srai x31 x31 3      ====        srai t6, t6, 3
                                                  30'd    6748    : data = 32'h    2B988113    ;    //    addi x2 x17 697      ====        addi sp, a7, 697
                                                  30'd    6749    : data = 32'h    00F49133    ;    //    sll x2 x9 x15      ====        sll sp, s1, a5
                                                  30'd    6750    : data = 32'h    00AEBE33    ;    //    sltu x28 x29 x10      ====        sltu t3, t4, a0
                                                  30'd    6751    : data = 32'h    41EBD813    ;    //    srai x16 x23 30      ====        srai a6, s7, 30
                                                  30'd    6752    : data = 32'h    3E2D9097    ;    //    auipc x1 254681      ====        auipc ra, 254681
                                                  30'd    6753    : data = 32'h    504E3C93    ;    //    sltiu x25 x28 1284      ====        sltiu s9, t3, 1284
                                                  30'd    6754    : data = 32'h    41408E33    ;    //    sub x28 x1 x20      ====        sub t3, ra, s4
                                                  30'd    6755    : data = 32'h    417888B3    ;    //    sub x17 x17 x23      ====        sub a7, a7, s7
                                                  30'd    6756    : data = 32'h    8AFC6B13    ;    //    ori x22 x24 -1873      ====        ori s6, s8, -1873
                                                  30'd    6757    : data = 32'h    00F8A1B3    ;    //    slt x3 x17 x15      ====        slt gp, a7, a5
                                                  30'd    6758    : data = 32'h    000D1333    ;    //    sll x6 x26 x0      ====        sll t1, s10, zero
                                                  30'd    6759    : data = 32'h    C861B713    ;    //    sltiu x14 x3 -890      ====        sltiu a4, gp, -890
                                                  30'd    6760    : data = 32'h    7AC85137    ;    //    lui x2 502917      ====        lui sp, 502917
                                                  30'd    6761    : data = 32'h    81E57117    ;    //    auipc x2 532055      ====        auipc sp, 532055
                                                  30'd    6762    : data = 32'h    01B6DA33    ;    //    srl x20 x13 x27      ====        srl s4, a3, s11
                                                  30'd    6763    : data = 32'h    01711733    ;    //    sll x14 x2 x23      ====        sll a4, sp, s7
                                                  30'd    6764    : data = 32'h    41A3D8B3    ;    //    sra x17 x7 x26      ====        sra a7, t2, s10
                                                  30'd    6765    : data = 32'h    01C75E33    ;    //    srl x28 x14 x28      ====        srl t3, a4, t3
                                                  30'd    6766    : data = 32'h    01F90433    ;    //    add x8 x18 x31      ====        add s0, s2, t6
                                                  30'd    6767    : data = 32'h    01905E33    ;    //    srl x28 x0 x25      ====        srl t3, zero, s9
                                                  30'd    6768    : data = 32'h    00EBCBB3    ;    //    xor x23 x23 x14      ====        xor s7, s7, a4
                                                  30'd    6769    : data = 32'h    ED30B793    ;    //    sltiu x15 x1 -301      ====        sltiu a5, ra, -301
                                                  30'd    6770    : data = 32'h    007FC733    ;    //    xor x14 x31 x7      ====        xor a4, t6, t2
                                                  30'd    6771    : data = 32'h    0196CEB3    ;    //    xor x29 x13 x25      ====        xor t4, a3, s9
                                                  30'd    6772    : data = 32'h    E980F0B7    ;    //    lui x1 956431      ====        lui ra, 956431
                                                  30'd    6773    : data = 32'h    01E6D7B3    ;    //    srl x15 x13 x30      ====        srl a5, a3, t5
                                                  30'd    6774    : data = 32'h    1B6EE097    ;    //    auipc x1 112366      ====        auipc ra, 112366
                                                  30'd    6775    : data = 32'h    0016D133    ;    //    srl x2 x13 x1      ====        srl sp, a3, ra
                                                  30'd    6776    : data = 32'h    017F1C93    ;    //    slli x25 x30 23      ====        slli s9, t5, 23
                                                  30'd    6777    : data = 32'h    C3076713    ;    //    ori x14 x14 -976      ====        ori a4, a4, -976
                                                  30'd    6778    : data = 32'h    005E9B13    ;    //    slli x22 x29 5      ====        slli s6, t4, 5
                                                  30'd    6779    : data = 32'h    3B786C13    ;    //    ori x24 x16 951      ====        ori s8, a6, 951
                                                  30'd    6780    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6781    : data = 32'h    01EFB0B3    ;    //    sltu x1 x31 x30      ====        sltu ra, t6, t5
                                                  30'd    6782    : data = 32'h    019D5E33    ;    //    srl x28 x26 x25      ====        srl t3, s10, s9
                                                  30'd    6783    : data = 32'h    2757E493    ;    //    ori x9 x15 629      ====        ori s1, a5, 629
                                                  30'd    6784    : data = 32'h    E9E14B93    ;    //    xori x23 x2 -354      ====        xori s7, sp, -354
                                                  30'd    6785    : data = 32'h    016C1333    ;    //    sll x6 x24 x22      ====        sll t1, s8, s6
                                                  30'd    6786    : data = 32'h    C7838913    ;    //    addi x18 x7 -904      ====        addi s2, t2, -904
                                                  30'd    6787    : data = 32'h    82624F93    ;    //    xori x31 x4 -2010      ====        xori t6, tp, -2010
                                                  30'd    6788    : data = 32'h    41D3DE13    ;    //    srai x28 x7 29      ====        srai t3, t2, 29
                                                  30'd    6789    : data = 32'h    019A1633    ;    //    sll x12 x20 x25      ====        sll a2, s4, s9
                                                  30'd    6790    : data = 32'h    C325C893    ;    //    xori x17 x11 -974      ====        xori a7, a1, -974
                                                  30'd    6791    : data = 32'h    EDCE6F93    ;    //    ori x31 x28 -292      ====        ori t6, t3, -292
                                                  30'd    6792    : data = 32'h    01EF0B33    ;    //    add x22 x30 x30      ====        add s6, t5, t5
                                                  30'd    6793    : data = 32'h    000D0933    ;    //    add x18 x26 x0      ====        add s2, s10, zero
                                                  30'd    6794    : data = 32'h    CAE3F993    ;    //    andi x19 x7 -850      ====        andi s3, t2, -850
                                                  30'd    6795    : data = 32'h    FFF00393    ;    //    addi x7 x0 -1      ====        li t2, 0xffffffff #start riscv_int_numeric_corner_stream_23
                                                  30'd    6796    : data = 32'h    733C2CB7    ;    //    lui x25 472002      ====        li s9, 0x733c21aa
                                                  30'd    6797    : data = 32'h    1AAC8C93    ;    //    addi x25 x25 426      ====        li s9, 0x733c21aa
                                                  30'd    6798    : data = 32'h    00000E13    ;    //    addi x28 x0 0      ====        li t3, 0x0
                                                  30'd    6799    : data = 32'h    80000637    ;    //    lui x12 524288      ====        li a2, 0x80000000
                                                  30'd    6800    : data = 32'h    00060613    ;    //    addi x12 x12 0      ====        li a2, 0x80000000
                                                  30'd    6801    : data = 32'h    F333DFB7    ;    //    lui x31 996157      ====        li t6, 0xf333d20b
                                                  30'd    6802    : data = 32'h    20BF8F93    ;    //    addi x31 x31 523      ====        li t6, 0xf333d20b
                                                  30'd    6803    : data = 32'h    FFF00A13    ;    //    addi x20 x0 -1      ====        li s4, 0xffffffff
                                                  30'd    6804    : data = 32'h    80000437    ;    //    lui x8 524288      ====        li s0, 0x80000000
                                                  30'd    6805    : data = 32'h    00040413    ;    //    addi x8 x8 0      ====        li s0, 0x80000000
                                                  30'd    6806    : data = 32'h    6CEF3837    ;    //    lui x16 446195      ====        li a6, 0x6cef2bf6
                                                  30'd    6807    : data = 32'h    BF680813    ;    //    addi x16 x16 -1034      ====        li a6, 0x6cef2bf6
                                                  30'd    6808    : data = 32'h    80000C37    ;    //    lui x24 524288      ====        li s8, 0x80000000
                                                  30'd    6809    : data = 32'h    000C0C13    ;    //    addi x24 x24 0      ====        li s8, 0x80000000
                                                  30'd    6810    : data = 32'h    FFF00693    ;    //    addi x13 x0 -1      ====        li a3, 0xffffffff
                                                  30'd    6811    : data = 32'h    00DC8CB3    ;    //    add x25 x25 x13      ====        add s9, s9, a3
                                                  30'd    6812    : data = 32'h    007E0FB3    ;    //    add x31 x28 x7      ====        add t6, t3, t2
                                                  30'd    6813    : data = 32'h    E5438693    ;    //    addi x13 x7 -428      ====        addi a3, t2, -428
                                                  30'd    6814    : data = 32'h    40D60A33    ;    //    sub x20 x12 x13      ====        sub s4, a2, a3
                                                  30'd    6815    : data = 32'h    41080833    ;    //    sub x16 x16 x16      ====        sub a6, a6, a6
                                                  30'd    6816    : data = 32'h    AC1C1A17    ;    //    auipc x20 704961      ====        auipc s4, 704961
                                                  30'd    6817    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6818    : data = 32'h    01C40FB3    ;    //    add x31 x8 x28      ====        add t6, s0, t3
                                                  30'd    6819    : data = 32'h    41C60A33    ;    //    sub x20 x12 x28      ====        sub s4, a2, t3
                                                  30'd    6820    : data = 32'h    008A0A33    ;    //    add x20 x20 x8      ====        add s4, s4, s0
                                                  30'd    6821    : data = 32'h    83F3CA17    ;    //    auipc x20 540476      ====        auipc s4, 540476
                                                  30'd    6822    : data = 32'h    AD02B3B7    ;    //    lui x7 708651      ====        lui t2, 708651
                                                  30'd    6823    : data = 32'h    40840C33    ;    //    sub x24 x8 x8      ====        sub s8, s0, s0
                                                  30'd    6824    : data = 32'h    AA6C8413    ;    //    addi x8 x25 -1370      ====        addi s0, s9, -1370
                                                  30'd    6825    : data = 32'h    268ADCB7    ;    //    lui x25 157869      ====        lui s9, 157869
                                                  30'd    6826    : data = 32'h    40C383B3    ;    //    sub x7 x7 x12      ====        sub t2, t2, a2
                                                  30'd    6827    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6828    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6829    : data = 32'h    435040EF    ;    //    jal x1 19508      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_23
                                                  30'd    6830    : data = 32'h    40645E13    ;    //    srai x28 x8 6      ====        srai t3, s0, 6
                                                  30'd    6831    : data = 32'h    011F1B93    ;    //    slli x23 x30 17      ====        slli s7, t5, 17
                                                  30'd    6832    : data = 32'h    16FED937    ;    //    lui x18 94189      ====        lui s2, 94189
                                                  30'd    6833    : data = 32'h    7FA94A93    ;    //    xori x21 x18 2042      ====        xori s5, s2, 2042
                                                  30'd    6834    : data = 32'h    408D81B3    ;    //    sub x3 x27 x8      ====        sub gp, s11, s0
                                                  30'd    6835    : data = 32'h    33C8A917    ;    //    auipc x18 212106      ====        auipc s2, 212106
                                                  30'd    6836    : data = 32'h    015BDA33    ;    //    srl x20 x23 x21      ====        srl s4, s7, s5
                                                  30'd    6837    : data = 32'h    F263E413    ;    //    ori x8 x7 -218      ====        ori s0, t2, -218
                                                  30'd    6838    : data = 32'h    01EE1933    ;    //    sll x18 x28 x30      ====        sll s2, t3, t5
                                                  30'd    6839    : data = 32'h    1A9D6493    ;    //    ori x9 x26 425      ====        ori s1, s10, 425
                                                  30'd    6840    : data = 32'h    006737B3    ;    //    sltu x15 x14 x6      ====        sltu a5, a4, t1
                                                  30'd    6841    : data = 32'h    01CCB297    ;    //    auipc x5 7371      ====        auipc t0, 7371
                                                  30'd    6842    : data = 32'h    011BB433    ;    //    sltu x8 x23 x17      ====        sltu s0, s7, a7
                                                  30'd    6843    : data = 32'h    01E81413    ;    //    slli x8 x16 30      ====        slli s0, a6, 30
                                                  30'd    6844    : data = 32'h    009DDE13    ;    //    srli x28 x27 9      ====        srli t3, s11, 9
                                                  30'd    6845    : data = 32'h    40E68D33    ;    //    sub x26 x13 x14      ====        sub s10, a3, a4
                                                  30'd    6846    : data = 32'h    005D5033    ;    //    srl x0 x26 x5      ====        srl zero, s10, t0
                                                  30'd    6847    : data = 32'h    853B0337    ;    //    lui x6 545712      ====        lui t1, 545712
                                                  30'd    6848    : data = 32'h    200C6E13    ;    //    ori x28 x24 512      ====        ori t3, s8, 512
                                                  30'd    6849    : data = 32'h    4019DD93    ;    //    srai x27 x19 1      ====        srai s11, s3, 1
                                                  30'd    6850    : data = 32'h    735B37B7    ;    //    lui x15 472499      ====        lui a5, 472499
                                                  30'd    6851    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6852    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6853    : data = 32'h    F70DCF93    ;    //    xori x31 x27 -144      ====        xori t6, s11, -144
                                                  30'd    6854    : data = 32'h    01A93E33    ;    //    sltu x28 x18 x26      ====        sltu t3, s2, s10
                                                  30'd    6855    : data = 32'h    411101B3    ;    //    sub x3 x2 x17      ====        sub gp, sp, a7
                                                  30'd    6856    : data = 32'h    87A7B613    ;    //    sltiu x12 x15 -1926      ====        sltiu a2, a5, -1926
                                                  30'd    6857    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6858    : data = 32'h    236DED93    ;    //    ori x27 x27 566      ====        ori s11, s11, 566
                                                  30'd    6859    : data = 32'h    016A9793    ;    //    slli x15 x21 22      ====        slli a5, s5, 22
                                                  30'd    6860    : data = 32'h    C8C58613    ;    //    addi x12 x11 -884      ====        addi a2, a1, -884
                                                  30'd    6861    : data = 32'h    00A31133    ;    //    sll x2 x6 x10      ====        sll sp, t1, a0
                                                  30'd    6862    : data = 32'h    DB173AB7    ;    //    lui x21 897395      ====        lui s5, 897395
                                                  30'd    6863    : data = 32'h    401CD0B3    ;    //    sra x1 x25 x1      ====        sra ra, s9, ra
                                                  30'd    6864    : data = 32'h    8550AF93    ;    //    slti x31 x1 -1963      ====        slti t6, ra, -1963
                                                  30'd    6865    : data = 32'h    DBB24D13    ;    //    xori x26 x4 -581      ====        xori s10, tp, -581
                                                  30'd    6866    : data = 32'h    00BDFB33    ;    //    and x22 x27 x11      ====        and s6, s11, a1
                                                  30'd    6867    : data = 32'h    4104D893    ;    //    srai x17 x9 16      ====        srai a7, s1, 16
                                                  30'd    6868    : data = 32'h    015D9633    ;    //    sll x12 x27 x21      ====        sll a2, s11, s5
                                                  30'd    6869    : data = 32'h    00A1BA33    ;    //    sltu x20 x3 x10      ====        sltu s4, gp, a0
                                                  30'd    6870    : data = 32'h    00B7ADB3    ;    //    slt x27 x15 x11      ====        slt s11, a5, a1
                                                  30'd    6871    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6872    : data = 32'h    01B1E033    ;    //    or x0 x3 x27      ====        or zero, gp, s11
                                                  30'd    6873    : data = 32'h    AB0C3593    ;    //    sltiu x11 x24 -1360      ====        sltiu a1, s8, -1360
                                                  30'd    6874    : data = 32'h    4047DA13    ;    //    srai x20 x15 4      ====        srai s4, a5, 4
                                                  30'd    6875    : data = 32'h    4B6B7493    ;    //    andi x9 x22 1206      ====        andi s1, s6, 1206
                                                  30'd    6876    : data = 32'h    014365B3    ;    //    or x11 x6 x20      ====        or a1, t1, s4
                                                  30'd    6877    : data = 32'h    C439C993    ;    //    xori x19 x19 -957      ====        xori s3, s3, -957
                                                  30'd    6878    : data = 32'h    68A02013    ;    //    slti x0 x0 1674      ====        slti zero, zero, 1674
                                                  30'd    6879    : data = 32'h    CFBC3037    ;    //    lui x0 850883      ====        lui zero, 850883
                                                  30'd    6880    : data = 32'h    66E9F113    ;    //    andi x2 x19 1646      ====        andi sp, s3, 1646
                                                  30'd    6881    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6882    : data = 32'h    40875433    ;    //    sra x8 x14 x8      ====        sra s0, a4, s0
                                                  30'd    6883    : data = 32'h    000B7833    ;    //    and x16 x22 x0      ====        and a6, s6, zero
                                                  30'd    6884    : data = 32'h    06262D17    ;    //    auipc x26 25186      ====        auipc s10, 25186
                                                  30'd    6885    : data = 32'h    0019D013    ;    //    srli x0 x19 1      ====        srli zero, s3, 1
                                                  30'd    6886    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6887    : data = 32'h    9146CA13    ;    //    xori x20 x13 -1772      ====        xori s4, a3, -1772
                                                  30'd    6888    : data = 32'h    024F4813    ;    //    xori x16 x30 36      ====        xori a6, t5, 36
                                                  30'd    6889    : data = 32'h    40AC5413    ;    //    srai x8 x24 10      ====        srai s0, s8, 10
                                                  30'd    6890    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6891    : data = 32'h    01DBCEB3    ;    //    xor x29 x23 x29      ====        xor t4, s7, t4
                                                  30'd    6892    : data = 32'h    00F80CB3    ;    //    add x25 x16 x15      ====        add s9, a6, a5
                                                  30'd    6893    : data = 32'h    AB5A45B7    ;    //    lui x11 701860      ====        lui a1, 701860
                                                  30'd    6894    : data = 32'h    00BE0E33    ;    //    add x28 x28 x11      ====        add t3, t3, a1
                                                  30'd    6895    : data = 32'h    38CCF013    ;    //    andi x0 x25 908      ====        andi zero, s9, 908
                                                  30'd    6896    : data = 32'h    406FD5B3    ;    //    sra x11 x31 x6      ====        sra a1, t6, t1
                                                  30'd    6897    : data = 32'h    FD260713    ;    //    addi x14 x12 -46      ====        addi a4, a2, -46
                                                  30'd    6898    : data = 32'h    E05264B7    ;    //    lui x9 918822      ====        lui s1, 918822
                                                  30'd    6899    : data = 32'h    000A0CB3    ;    //    add x25 x20 x0      ====        add s9, s4, zero
                                                  30'd    6900    : data = 32'h    00EAAA33    ;    //    slt x20 x21 x14      ====        slt s4, s5, a4
                                                  30'd    6901    : data = 32'h    00968633    ;    //    add x12 x13 x9      ====        add a2, a3, s1
                                                  30'd    6902    : data = 32'h    F7152913    ;    //    slti x18 x10 -143      ====        slti s2, a0, -143
                                                  30'd    6903    : data = 32'h    00FD1AB3    ;    //    sll x21 x26 x15      ====        sll s5, s10, a5
                                                  30'd    6904    : data = 32'h    0080A0B3    ;    //    slt x1 x1 x8      ====        slt ra, ra, s0
                                                  30'd    6905    : data = 32'h    013484B3    ;    //    add x9 x9 x19      ====        add s1, s1, s3
                                                  30'd    6906    : data = 32'h    7CC50013    ;    //    addi x0 x10 1996      ====        addi zero, a0, 1996
                                                  30'd    6907    : data = 32'h    D59DCE93    ;    //    xori x29 x27 -679      ====        xori t4, s11, -679
                                                  30'd    6908    : data = 32'h    011E1893    ;    //    slli x17 x28 17      ====        slli a7, t3, 17
                                                  30'd    6909    : data = 32'h    D28F2613    ;    //    slti x12 x30 -728      ====        slti a2, t5, -728
                                                  30'd    6910    : data = 32'h    00B54CB3    ;    //    xor x25 x10 x11      ====        xor s9, a0, a1
                                                  30'd    6911    : data = 32'h    00517E33    ;    //    and x28 x2 x5      ====        and t3, sp, t0
                                                  30'd    6912    : data = 32'h    2D5EFF93    ;    //    andi x31 x29 725      ====        andi t6, t4, 725
                                                  30'd    6913    : data = 32'h    00BC1093    ;    //    slli x1 x24 11      ====        slli ra, s8, 11
                                                  30'd    6914    : data = 32'h    00F2DF93    ;    //    srli x31 x5 15      ====        srli t6, t0, 15
                                                  30'd    6915    : data = 32'h    00551F93    ;    //    slli x31 x10 5      ====        slli t6, a0, 5
                                                  30'd    6916    : data = 32'h    4131D913    ;    //    srai x18 x3 19      ====        srai s2, gp, 19
                                                  30'd    6917    : data = 32'h    01BDFEB3    ;    //    and x29 x27 x27      ====        and t4, s11, s11
                                                  30'd    6918    : data = 32'h    00C545B3    ;    //    xor x11 x10 x12      ====        xor a1, a0, a2
                                                  30'd    6919    : data = 32'h    44108013    ;    //    addi x0 x1 1089      ====        addi zero, ra, 1089
                                                  30'd    6920    : data = 32'h    A41A3D93    ;    //    sltiu x27 x20 -1471      ====        sltiu s11, s4, -1471
                                                  30'd    6921    : data = 32'h    7F0D6293    ;    //    ori x5 x26 2032      ====        ori t0, s10, 2032
                                                  30'd    6922    : data = 32'h    C647A093    ;    //    slti x1 x15 -924      ====        slti ra, a5, -924
                                                  30'd    6923    : data = 32'h    9211E913    ;    //    ori x18 x3 -1759      ====        ori s2, gp, -1759
                                                  30'd    6924    : data = 32'h    6CBA42B7    ;    //    lui x5 445348      ====        lui t0, 445348
                                                  30'd    6925    : data = 32'h    41ECD893    ;    //    srai x17 x25 30      ====        srai a7, s9, 30
                                                  30'd    6926    : data = 32'h    1DC54593    ;    //    xori x11 x10 476      ====        xori a1, a0, 476
                                                  30'd    6927    : data = 32'h    BFFBEB13    ;    //    ori x22 x23 -1025      ====        ori s6, s7, -1025
                                                  30'd    6928    : data = 32'h    E27D4E93    ;    //    xori x29 x26 -473      ====        xori t4, s10, -473
                                                  30'd    6929    : data = 32'h    00A2CFB3    ;    //    xor x31 x5 x10      ====        xor t6, t0, a0
                                                  30'd    6930    : data = 32'h    003607B3    ;    //    add x15 x12 x3      ====        add a5, a2, gp
                                                  30'd    6931    : data = 32'h    41D58D33    ;    //    sub x26 x11 x29      ====        sub s10, a1, t4
                                                  30'd    6932    : data = 32'h    014676B3    ;    //    and x13 x12 x20      ====        and a3, a2, s4
                                                  30'd    6933    : data = 32'h    00A96B33    ;    //    or x22 x18 x10      ====        or s6, s2, a0
                                                  30'd    6934    : data = 32'h    4B696013    ;    //    ori x0 x18 1206      ====        ori zero, s2, 1206
                                                  30'd    6935    : data = 32'h    00FE73B3    ;    //    and x7 x28 x15      ====        and t2, t3, a5
                                                  30'd    6936    : data = 32'h    00491BB3    ;    //    sll x23 x18 x4      ====        sll s7, s2, tp
                                                  30'd    6937    : data = 32'h    9B437013    ;    //    andi x0 x6 -1612      ====        andi zero, t1, -1612
                                                  30'd    6938    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6939    : data = 32'h    002D40B3    ;    //    xor x1 x26 x2      ====        xor ra, s10, sp
                                                  30'd    6940    : data = 32'h    F600CC13    ;    //    xori x24 x1 -160      ====        xori s8, ra, -160
                                                  30'd    6941    : data = 32'h    CAF58793    ;    //    addi x15 x11 -849      ====        addi a5, a1, -849
                                                  30'd    6942    : data = 32'h    00591E33    ;    //    sll x28 x18 x5      ====        sll t3, s2, t0
                                                  30'd    6943    : data = 32'h    01C367B3    ;    //    or x15 x6 x28      ====        or a5, t1, t3
                                                  30'd    6944    : data = 32'h    00C77A33    ;    //    and x20 x14 x12      ====        and s4, a4, a2
                                                  30'd    6945    : data = 32'h    21A5AD93    ;    //    slti x27 x11 538      ====        slti s11, a1, 538
                                                  30'd    6946    : data = 32'h    0043F2B3    ;    //    and x5 x7 x4      ====        and t0, t2, tp
                                                  30'd    6947    : data = 32'h    5D70CA93    ;    //    xori x21 x1 1495      ====        xori s5, ra, 1495
                                                  30'd    6948    : data = 32'h    5D000DB7    ;    //    lui x27 380928      ====        lui s11, 380928
                                                  30'd    6949    : data = 32'h    01654A33    ;    //    xor x20 x10 x22      ====        xor s4, a0, s6
                                                  30'd    6950    : data = 32'h    015BF5B3    ;    //    and x11 x23 x21      ====        and a1, s7, s5
                                                  30'd    6951    : data = 32'h    00EA9593    ;    //    slli x11 x21 14      ====        slli a1, s5, 14
                                                  30'd    6952    : data = 32'h    015ABA13    ;    //    sltiu x20 x21 21      ====        sltiu s4, s5, 21
                                                  30'd    6953    : data = 32'h    8F36C393    ;    //    xori x7 x13 -1805      ====        xori t2, a3, -1805
                                                  30'd    6954    : data = 32'h    00462933    ;    //    slt x18 x12 x4      ====        slt s2, a2, tp
                                                  30'd    6955    : data = 32'h    00429BB3    ;    //    sll x23 x5 x4      ====        sll s7, t0, tp
                                                  30'd    6956    : data = 32'h    AEEE8297    ;    //    auipc x5 716520      ====        auipc t0, 716520
                                                  30'd    6957    : data = 32'h    00B75D93    ;    //    srli x27 x14 11      ====        srli s11, a4, 11
                                                  30'd    6958    : data = 32'h    0180A733    ;    //    slt x14 x1 x24      ====        slt a4, ra, s8
                                                  30'd    6959    : data = 32'h    011FBFB3    ;    //    sltu x31 x31 x17      ====        sltu t6, t6, a7
                                                  30'd    6960    : data = 32'h    0170EBB3    ;    //    or x23 x1 x23      ====        or s7, ra, s7
                                                  30'd    6961    : data = 32'h    59183093    ;    //    sltiu x1 x16 1425      ====        sltiu ra, a6, 1425
                                                  30'd    6962    : data = 32'h    D09C36B7    ;    //    lui x13 854467      ====        lui a3, 854467
                                                  30'd    6963    : data = 32'h    015D8BB3    ;    //    add x23 x27 x21      ====        add s7, s11, s5
                                                  30'd    6964    : data = 32'h    005732B3    ;    //    sltu x5 x14 x5      ====        sltu t0, a4, t0
                                                  30'd    6965    : data = 32'h    B2EB6493    ;    //    ori x9 x22 -1234      ====        ori s1, s6, -1234
                                                  30'd    6966    : data = 32'h    00A682B3    ;    //    add x5 x13 x10      ====        add t0, a3, a0
                                                  30'd    6967    : data = 32'h    DE343A13    ;    //    sltiu x20 x8 -541      ====        sltiu s4, s0, -541
                                                  30'd    6968    : data = 32'h    DA3BD4B7    ;    //    lui x9 893885      ====        lui s1, 893885
                                                  30'd    6969    : data = 32'h    959E0D93    ;    //    addi x27 x28 -1703      ====        addi s11, t3, -1703
                                                  30'd    6970    : data = 32'h    002C1133    ;    //    sll x2 x24 x2      ====        sll sp, s8, sp
                                                  30'd    6971    : data = 32'h    41078D33    ;    //    sub x26 x15 x16      ====        sub s10, a5, a6
                                                  30'd    6972    : data = 32'h    0102F7B3    ;    //    and x15 x5 x16      ====        and a5, t0, a6
                                                  30'd    6973    : data = 32'h    FCDAF793    ;    //    andi x15 x21 -51      ====        andi a5, s5, -51
                                                  30'd    6974    : data = 32'h    00B765B3    ;    //    or x11 x14 x11      ====        or a1, a4, a1
                                                  30'd    6975    : data = 32'h    51714613    ;    //    xori x12 x2 1303      ====        xori a2, sp, 1303
                                                  30'd    6976    : data = 32'h    01261933    ;    //    sll x18 x12 x18      ====        sll s2, a2, s2
                                                  30'd    6977    : data = 32'h    01AD1313    ;    //    slli x6 x26 26      ====        slli t1, s10, 26
                                                  30'd    6978    : data = 32'h    F58AA813    ;    //    slti x16 x21 -168      ====        slti a6, s5, -168
                                                  30'd    6979    : data = 32'h    00C9E433    ;    //    or x8 x19 x12      ====        or s0, s3, a2
                                                  30'd    6980    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    6981    : data = 32'h    00D76DB3    ;    //    or x27 x14 x13      ====        or s11, a4, a3
                                                  30'd    6982    : data = 32'h    28BF6293    ;    //    ori x5 x30 651      ====        ori t0, t5, 651
                                                  30'd    6983    : data = 32'h    008BC4B3    ;    //    xor x9 x23 x8      ====        xor s1, s7, s0
                                                  30'd    6984    : data = 32'h    00152133    ;    //    slt x2 x10 x1      ====        slt sp, a0, ra
                                                  30'd    6985    : data = 32'h    010A6333    ;    //    or x6 x20 x16      ====        or t1, s4, a6
                                                  30'd    6986    : data = 32'h    0186D633    ;    //    srl x12 x13 x24      ====        srl a2, a3, s8
                                                  30'd    6987    : data = 32'h    00191833    ;    //    sll x16 x18 x1      ====        sll a6, s2, ra
                                                  30'd    6988    : data = 32'h    019D0E33    ;    //    add x28 x26 x25      ====        add t3, s10, s9
                                                  30'd    6989    : data = 32'h    01BC5833    ;    //    srl x16 x24 x27      ====        srl a6, s8, s11
                                                  30'd    6990    : data = 32'h    7FF52A13    ;    //    slti x20 x10 2047      ====        slti s4, a0, 2047
                                                  30'd    6991    : data = 32'h    B3514497    ;    //    auipc x9 734484      ====        auipc s1, 734484
                                                  30'd    6992    : data = 32'h    416609B3    ;    //    sub x19 x12 x22      ====        sub s3, a2, s6
                                                  30'd    6993    : data = 32'h    4140DD13    ;    //    srai x26 x1 20      ====        srai s10, ra, 20
                                                  30'd    6994    : data = 32'h    000ED1B3    ;    //    srl x3 x29 x0      ====        srl gp, t4, zero
                                                  30'd    6995    : data = 32'h    009E15B3    ;    //    sll x11 x28 x9      ====        sll a1, t3, s1
                                                  30'd    6996    : data = 32'h    00A8F633    ;    //    and x12 x17 x10      ====        and a2, a7, a0
                                                  30'd    6997    : data = 32'h    00FFCB33    ;    //    xor x22 x31 x15      ====        xor s6, t6, a5
                                                  30'd    6998    : data = 32'h    B5849317    ;    //    auipc x6 743497      ====        auipc t1, 743497
                                                  30'd    6999    : data = 32'h    CDA3BD13    ;    //    sltiu x26 x7 -806      ====        sltiu s10, t2, -806
                                                  30'd    7000    : data = 32'h    26184293    ;    //    xori x5 x16 609      ====        xori t0, a6, 609
                                                  30'd    7001    : data = 32'h    01DAF4B3    ;    //    and x9 x21 x29      ====        and s1, s5, t4
                                                  30'd    7002    : data = 32'h    F806AE93    ;    //    slti x29 x13 -128      ====        slti t4, a3, -128
                                                  30'd    7003    : data = 32'h    62A8C613    ;    //    xori x12 x17 1578      ====        xori a2, a7, 1578
                                                  30'd    7004    : data = 32'h    CAF0C413    ;    //    xori x8 x1 -849      ====        xori s0, ra, -849
                                                  30'd    7005    : data = 32'h    D8726693    ;    //    ori x13 x4 -633      ====        ori a3, tp, -633
                                                  30'd    7006    : data = 32'h    00825293    ;    //    srli x5 x4 8      ====        srli t0, tp, 8
                                                  30'd    7007    : data = 32'h    BD66B817    ;    //    auipc x16 775787      ====        auipc a6, 775787
                                                  30'd    7008    : data = 32'h    3EB56893    ;    //    ori x17 x10 1003      ====        ori a7, a0, 1003
                                                  30'd    7009    : data = 32'h    65CEB117    ;    //    auipc x2 417003      ====        auipc sp, 417003
                                                  30'd    7010    : data = 32'h    01F59913    ;    //    slli x18 x11 31      ====        slli s2, a1, 31
                                                  30'd    7011    : data = 32'h    8339E613    ;    //    ori x12 x19 -1997      ====        ori a2, s3, -1997
                                                  30'd    7012    : data = 32'h    FB3924B7    ;    //    lui x9 1029010      ====        lui s1, 1029010
                                                  30'd    7013    : data = 32'h    F235B993    ;    //    sltiu x19 x11 -221      ====        sltiu s3, a1, -221
                                                  30'd    7014    : data = 32'h    00B948B3    ;    //    xor x17 x18 x11      ====        xor a7, s2, a1
                                                  30'd    7015    : data = 32'h    012AEE33    ;    //    or x28 x21 x18      ====        or t3, s5, s2
                                                  30'd    7016    : data = 32'h    4CC06E13    ;    //    ori x28 x0 1228      ====        ori t3, zero, 1228
                                                  30'd    7017    : data = 32'h    40755B13    ;    //    srai x22 x10 7      ====        srai s6, a0, 7
                                                  30'd    7018    : data = 32'h    5C373693    ;    //    sltiu x13 x14 1475      ====        sltiu a3, a4, 1475
                                                  30'd    7019    : data = 32'h    00406733    ;    //    or x14 x0 x4      ====        or a4, zero, tp
                                                  30'd    7020    : data = 32'h    01BE1B13    ;    //    slli x22 x28 27      ====        slli s6, t3, 27
                                                  30'd    7021    : data = 32'h    004BBAB3    ;    //    sltu x21 x23 x4      ====        sltu s5, s7, tp
                                                  30'd    7022    : data = 32'h    01D576B3    ;    //    and x13 x10 x29      ====        and a3, a0, t4
                                                  30'd    7023    : data = 32'h    FAB6B593    ;    //    sltiu x11 x13 -85      ====        sltiu a1, a3, -85
                                                  30'd    7024    : data = 32'h    37543737    ;    //    lui x14 226627      ====        lui a4, 226627
                                                  30'd    7025    : data = 32'h    01E5DDB3    ;    //    srl x27 x11 x30      ====        srl s11, a1, t5
                                                  30'd    7026    : data = 32'h    015832B3    ;    //    sltu x5 x16 x21      ====        sltu t0, a6, s5
                                                  30'd    7027    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7028    : data = 32'h    7633FF93    ;    //    andi x31 x7 1891      ====        andi t6, t2, 1891
                                                  30'd    7029    : data = 32'h    6E637E13    ;    //    andi x28 x6 1766      ====        andi t3, t1, 1766
                                                  30'd    7030    : data = 32'h    37503B93    ;    //    sltiu x23 x0 885      ====        sltiu s7, zero, 885
                                                  30'd    7031    : data = 32'h    ECE18693    ;    //    addi x13 x3 -306      ====        addi a3, gp, -306
                                                  30'd    7032    : data = 32'h    FB104793    ;    //    xori x15 x0 -79      ====        xori a5, zero, -79
                                                  30'd    7033    : data = 32'h    72D14837    ;    //    lui x16 470292      ====        lui a6, 470292
                                                  30'd    7034    : data = 32'h    00CBD313    ;    //    srli x6 x23 12      ====        srli t1, s7, 12
                                                  30'd    7035    : data = 32'h    4079DB13    ;    //    srai x22 x19 7      ====        srai s6, s3, 7
                                                  30'd    7036    : data = 32'h    000000B3    ;    //    add x1 x0 x0      ====        add ra, zero, zero
                                                  30'd    7037    : data = 32'h    01927333    ;    //    and x6 x4 x25      ====        and t1, tp, s9
                                                  30'd    7038    : data = 32'h    005ADA13    ;    //    srli x20 x21 5      ====        srli s4, s5, 5
                                                  30'd    7039    : data = 32'h    EE60B193    ;    //    sltiu x3 x1 -282      ====        sltiu gp, ra, -282
                                                  30'd    7040    : data = 32'h    00C57733    ;    //    and x14 x10 x12      ====        and a4, a0, a2
                                                  30'd    7041    : data = 32'h    012559B3    ;    //    srl x19 x10 x18      ====        srl s3, a0, s2
                                                  30'd    7042    : data = 32'h    D15AF693    ;    //    andi x13 x21 -747      ====        andi a3, s5, -747
                                                  30'd    7043    : data = 32'h    017C5333    ;    //    srl x6 x24 x23      ====        srl t1, s8, s7
                                                  30'd    7044    : data = 32'h    C4B80337    ;    //    lui x6 805760      ====        lui t1, 805760
                                                  30'd    7045    : data = 32'h    01E12AB3    ;    //    slt x21 x2 x30      ====        slt s5, sp, t5
                                                  30'd    7046    : data = 32'h    41855B33    ;    //    sra x22 x10 x24      ====        sra s6, a0, s8
                                                  30'd    7047    : data = 32'h    FCD64713    ;    //    xori x14 x12 -51      ====        xori a4, a2, -51
                                                  30'd    7048    : data = 32'h    CE3E2613    ;    //    slti x12 x28 -797      ====        slti a2, t3, -797
                                                  30'd    7049    : data = 32'h    017D2A33    ;    //    slt x20 x26 x23      ====        slt s4, s10, s7
                                                  30'd    7050    : data = 32'h    00C29333    ;    //    sll x6 x5 x12      ====        sll t1, t0, a2
                                                  30'd    7051    : data = 32'h    401D8333    ;    //    sub x6 x27 x1      ====        sub t1, s11, ra
                                                  30'd    7052    : data = 32'h    01339F93    ;    //    slli x31 x7 19      ====        slli t6, t2, 19
                                                  30'd    7053    : data = 32'h    37D88D13    ;    //    addi x26 x17 893      ====        addi s10, a7, 893
                                                  30'd    7054    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7055    : data = 32'h    1E664FB7    ;    //    lui x31 124516      ====        lui t6, 124516
                                                  30'd    7056    : data = 32'h    40920933    ;    //    sub x18 x4 x9      ====        sub s2, tp, s1
                                                  30'd    7057    : data = 32'h    006D6133    ;    //    or x2 x26 x6      ====        or sp, s10, t1
                                                  30'd    7058    : data = 32'h    CC292113    ;    //    slti x2 x18 -830      ====        slti sp, s2, -830
                                                  30'd    7059    : data = 32'h    00319DB3    ;    //    sll x27 x3 x3      ====        sll s11, gp, gp
                                                  30'd    7060    : data = 32'h    00CB29B3    ;    //    slt x19 x22 x12      ====        slt s3, s6, a2
                                                  30'd    7061    : data = 32'h    018A9B33    ;    //    sll x22 x21 x24      ====        sll s6, s5, s8
                                                  30'd    7062    : data = 32'h    015584B3    ;    //    add x9 x11 x21      ====        add s1, a1, s5
                                                  30'd    7063    : data = 32'h    00F7D9B3    ;    //    srl x19 x15 x15      ====        srl s3, a5, a5
                                                  30'd    7064    : data = 32'h    016A9F93    ;    //    slli x31 x21 22      ====        slli t6, s5, 22
                                                  30'd    7065    : data = 32'h    C8980793    ;    //    addi x15 x16 -887      ====        addi a5, a6, -887
                                                  30'd    7066    : data = 32'h    0194DD33    ;    //    srl x26 x9 x25      ====        srl s10, s1, s9
                                                  30'd    7067    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7068    : data = 32'h    40A7D8B3    ;    //    sra x17 x15 x10      ====        sra a7, a5, a0
                                                  30'd    7069    : data = 32'h    012E5E13    ;    //    srli x28 x28 18      ====        srli t3, t3, 18
                                                  30'd    7070    : data = 32'h    00ABC633    ;    //    xor x12 x23 x10      ====        xor a2, s7, a0
                                                  30'd    7071    : data = 32'h    004C8733    ;    //    add x14 x25 x4      ====        add a4, s9, tp
                                                  30'd    7072    : data = 32'h    00EB5EB3    ;    //    srl x29 x22 x14      ====        srl t4, s6, a4
                                                  30'd    7073    : data = 32'h    E964B913    ;    //    sltiu x18 x9 -362      ====        sltiu s2, s1, -362
                                                  30'd    7074    : data = 32'h    00110BB3    ;    //    add x23 x2 x1      ====        add s7, sp, ra
                                                  30'd    7075    : data = 32'h    D0657117    ;    //    auipc x2 853591      ====        auipc sp, 853591
                                                  30'd    7076    : data = 32'h    01CEDE33    ;    //    srl x28 x29 x28      ====        srl t3, t4, t3
                                                  30'd    7077    : data = 32'h    225DB293    ;    //    sltiu x5 x27 549      ====        sltiu t0, s11, 549
                                                  30'd    7078    : data = 32'h    0184DEB3    ;    //    srl x29 x9 x24      ====        srl t4, s1, s8
                                                  30'd    7079    : data = 32'h    018CC633    ;    //    xor x12 x25 x24      ====        xor a2, s9, s8
                                                  30'd    7080    : data = 32'h    01A5FAB3    ;    //    and x21 x11 x26      ====        and s5, a1, s10
                                                  30'd    7081    : data = 32'h    361BE413    ;    //    ori x8 x23 865      ====        ori s0, s7, 865
                                                  30'd    7082    : data = 32'h    011A5FB3    ;    //    srl x31 x20 x17      ====        srl t6, s4, a7
                                                  30'd    7083    : data = 32'h    01169FB3    ;    //    sll x31 x13 x17      ====        sll t6, a3, a7
                                                  30'd    7084    : data = 32'h    00491413    ;    //    slli x8 x18 4      ====        slli s0, s2, 4
                                                  30'd    7085    : data = 32'h    00CC7433    ;    //    and x8 x24 x12      ====        and s0, s8, a2
                                                  30'd    7086    : data = 32'h    DD2D3B13    ;    //    sltiu x22 x26 -558      ====        sltiu s6, s10, -558
                                                  30'd    7087    : data = 32'h    01359D93    ;    //    slli x27 x11 19      ====        slli s11, a1, 19
                                                  30'd    7088    : data = 32'h    4001DF93    ;    //    srai x31 x3 0      ====        srai t6, gp, 0
                                                  30'd    7089    : data = 32'h    01DF1BB3    ;    //    sll x23 x30 x29      ====        sll s7, t5, t4
                                                  30'd    7090    : data = 32'h    41DD0BB3    ;    //    sub x23 x26 x29      ====        sub s7, s10, t4
                                                  30'd    7091    : data = 32'h    2779E693    ;    //    ori x13 x19 631      ====        ori a3, s3, 631
                                                  30'd    7092    : data = 32'h    01A79833    ;    //    sll x16 x15 x26      ====        sll a6, a5, s10
                                                  30'd    7093    : data = 32'h    01B1F433    ;    //    and x8 x3 x27      ====        and s0, gp, s11
                                                  30'd    7094    : data = 32'h    A168B293    ;    //    sltiu x5 x17 -1514      ====        sltiu t0, a7, -1514
                                                  30'd    7095    : data = 32'h    01E51733    ;    //    sll x14 x10 x30      ====        sll a4, a0, t5
                                                  30'd    7096    : data = 32'h    40DF5793    ;    //    srai x15 x30 13      ====        srai a5, t5, 13
                                                  30'd    7097    : data = 32'h    0140B733    ;    //    sltu x14 x1 x20      ====        sltu a4, ra, s4
                                                  30'd    7098    : data = 32'h    E959C893    ;    //    xori x17 x19 -363      ====        xori a7, s3, -363
                                                  30'd    7099    : data = 32'h    D8527993    ;    //    andi x19 x4 -635      ====        andi s3, tp, -635
                                                  30'd    7100    : data = 32'h    3BCE6613    ;    //    ori x12 x28 956      ====        ori a2, t3, 956
                                                  30'd    7101    : data = 32'h    0053B8B3    ;    //    sltu x17 x7 x5      ====        sltu a7, t2, t0
                                                  30'd    7102    : data = 32'h    417FD333    ;    //    sra x6 x31 x23      ====        sra t1, t6, s7
                                                  30'd    7103    : data = 32'h    33633C13    ;    //    sltiu x24 x6 822      ====        sltiu s8, t1, 822
                                                  30'd    7104    : data = 32'h    01EDD493    ;    //    srli x9 x27 30      ====        srli s1, s11, 30
                                                  30'd    7105    : data = 32'h    E50C6A97    ;    //    auipc x21 938182      ====        auipc s5, 938182
                                                  30'd    7106    : data = 32'h    0DB60593    ;    //    addi x11 x12 219      ====        addi a1, a2, 219
                                                  30'd    7107    : data = 32'h    00ECE3B3    ;    //    or x7 x25 x14      ====        or t2, s9, a4
                                                  30'd    7108    : data = 32'h    00C6FEB3    ;    //    and x29 x13 x12      ====        and t4, a3, a2
                                                  30'd    7109    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7110    : data = 32'h    41D55D93    ;    //    srai x27 x10 29      ====        srai s11, a0, 29
                                                  30'd    7111    : data = 32'h    010263B3    ;    //    or x7 x4 x16      ====        or t2, tp, a6
                                                  30'd    7112    : data = 32'h    013E9B13    ;    //    slli x22 x29 19      ====        slli s6, t4, 19
                                                  30'd    7113    : data = 32'h    01D3A933    ;    //    slt x18 x7 x29      ====        slt s2, t2, t4
                                                  30'd    7114    : data = 32'h    01B53D33    ;    //    sltu x26 x10 x27      ====        sltu s10, a0, s11
                                                  30'd    7115    : data = 32'h    01E5D893    ;    //    srli x17 x11 30      ====        srli a7, a1, 30
                                                  30'd    7116    : data = 32'h    01769993    ;    //    slli x19 x13 23      ====        slli s3, a3, 23
                                                  30'd    7117    : data = 32'h    417951B3    ;    //    sra x3 x18 x23      ====        sra gp, s2, s7
                                                  30'd    7118    : data = 32'h    0082B193    ;    //    sltiu x3 x5 8      ====        sltiu gp, t0, 8
                                                  30'd    7119    : data = 32'h    01399993    ;    //    slli x19 x19 19      ====        slli s3, s3, 19
                                                  30'd    7120    : data = 32'h    404CD313    ;    //    srai x6 x25 4      ====        srai t1, s9, 4
                                                  30'd    7121    : data = 32'h    00F78DB3    ;    //    add x27 x15 x15      ====        add s11, a5, a5
                                                  30'd    7122    : data = 32'h    016DA833    ;    //    slt x16 x27 x22      ====        slt a6, s11, s6
                                                  30'd    7123    : data = 32'h    00B0D133    ;    //    srl x2 x1 x11      ====        srl sp, ra, a1
                                                  30'd    7124    : data = 32'h    00AE7A33    ;    //    and x20 x28 x10      ====        and s4, t3, a0
                                                  30'd    7125    : data = 32'h    411D59B3    ;    //    sra x19 x26 x17      ====        sra s3, s10, a7
                                                  30'd    7126    : data = 32'h    0003B633    ;    //    sltu x12 x7 x0      ====        sltu a2, t2, zero
                                                  30'd    7127    : data = 32'h    402ADF93    ;    //    srai x31 x21 2      ====        srai t6, s5, 2
                                                  30'd    7128    : data = 32'h    017E5033    ;    //    srl x0 x28 x23      ====        srl zero, t3, s7
                                                  30'd    7129    : data = 32'h    01485613    ;    //    srli x12 x16 20      ====        srli a2, a6, 20
                                                  30'd    7130    : data = 32'h    00BB8033    ;    //    add x0 x23 x11      ====        add zero, s7, a1
                                                  30'd    7131    : data = 32'h    D835E813    ;    //    ori x16 x11 -637      ====        ori a6, a1, -637
                                                  30'd    7132    : data = 32'h    292BF593    ;    //    andi x11 x23 658      ====        andi a1, s7, 658
                                                  30'd    7133    : data = 32'h    7782EB17    ;    //    auipc x22 489518      ====        auipc s6, 489518
                                                  30'd    7134    : data = 32'h    00C29193    ;    //    slli x3 x5 12      ====        slli gp, t0, 12
                                                  30'd    7135    : data = 32'h    69A8B393    ;    //    sltiu x7 x17 1690      ====        sltiu t2, a7, 1690
                                                  30'd    7136    : data = 32'h    91FD0E13    ;    //    addi x28 x26 -1761      ====        addi t3, s10, -1761
                                                  30'd    7137    : data = 32'h    41875733    ;    //    sra x14 x14 x24      ====        sra a4, a4, s8
                                                  30'd    7138    : data = 32'h    00A418B3    ;    //    sll x17 x8 x10      ====        sll a7, s0, a0
                                                  30'd    7139    : data = 32'h    00981693    ;    //    slli x13 x16 9      ====        slli a3, a6, 9
                                                  30'd    7140    : data = 32'h    27BA2793    ;    //    slti x15 x20 635      ====        slti a5, s4, 635
                                                  30'd    7141    : data = 32'h    01B1E933    ;    //    or x18 x3 x27      ====        or s2, gp, s11
                                                  30'd    7142    : data = 32'h    018457B3    ;    //    srl x15 x8 x24      ====        srl a5, s0, s8
                                                  30'd    7143    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7144    : data = 32'h    FFC49E97    ;    //    auipc x29 1047625      ====        auipc t4, 1047625
                                                  30'd    7145    : data = 32'h    012C71B3    ;    //    and x3 x24 x18      ====        and gp, s8, s2
                                                  30'd    7146    : data = 32'h    41690633    ;    //    sub x12 x18 x22      ====        sub a2, s2, s6
                                                  30'd    7147    : data = 32'h    005072B3    ;    //    and x5 x0 x5      ====        and t0, zero, t0
                                                  30'd    7148    : data = 32'h    00AFC7B3    ;    //    xor x15 x31 x10      ====        xor a5, t6, a0
                                                  30'd    7149    : data = 32'h    0198D593    ;    //    srli x11 x17 25      ====        srli a1, a7, 25
                                                  30'd    7150    : data = 32'h    01EE71B3    ;    //    and x3 x28 x30      ====        and gp, t3, t5
                                                  30'd    7151    : data = 32'h    3E61AA13    ;    //    slti x20 x3 998      ====        slti s4, gp, 998
                                                  30'd    7152    : data = 32'h    008B5FB3    ;    //    srl x31 x22 x8      ====        srl t6, s6, s0
                                                  30'd    7153    : data = 32'h    007482B3    ;    //    add x5 x9 x7      ====        add t0, s1, t2
                                                  30'd    7154    : data = 32'h    01D3CC33    ;    //    xor x24 x7 x29      ====        xor s8, t2, t4
                                                  30'd    7155    : data = 32'h    B03B8637    ;    //    lui x12 721848      ====        lui a2, 721848
                                                  30'd    7156    : data = 32'h    002D8DB3    ;    //    add x27 x27 x2      ====        add s11, s11, sp
                                                  30'd    7157    : data = 32'h    01DB5713    ;    //    srli x14 x22 29      ====        srli a4, s6, 29
                                                  30'd    7158    : data = 32'h    00A1BEB3    ;    //    sltu x29 x3 x10      ====        sltu t4, gp, a0
                                                  30'd    7159    : data = 32'h    00B4D433    ;    //    srl x8 x9 x11      ====        srl s0, s1, a1
                                                  30'd    7160    : data = 32'h    00B331B3    ;    //    sltu x3 x6 x11      ====        sltu gp, t1, a1
                                                  30'd    7161    : data = 32'h    009D1B13    ;    //    slli x22 x26 9      ====        slli s6, s10, 9
                                                  30'd    7162    : data = 32'h    003835B3    ;    //    sltu x11 x16 x3      ====        sltu a1, a6, gp
                                                  30'd    7163    : data = 32'h    003FADB3    ;    //    slt x27 x31 x3      ====        slt s11, t6, gp
                                                  30'd    7164    : data = 32'h    00552733    ;    //    slt x14 x10 x5      ====        slt a4, a0, t0
                                                  30'd    7165    : data = 32'h    0EE6FC93    ;    //    andi x25 x13 238      ====        andi s9, a3, 238
                                                  30'd    7166    : data = 32'h    9B394A93    ;    //    xori x21 x18 -1613      ====        xori s5, s2, -1613
                                                  30'd    7167    : data = 32'h    41068B33    ;    //    sub x22 x13 x16      ====        sub s6, a3, a6
                                                  30'd    7168    : data = 32'h    016F1293    ;    //    slli x5 x30 22      ====        slli t0, t5, 22
                                                  30'd    7169    : data = 32'h    00FE1C93    ;    //    slli x25 x28 15      ====        slli s9, t3, 15
                                                  30'd    7170    : data = 32'h    4689FD93    ;    //    andi x27 x19 1128      ====        andi s11, s3, 1128
                                                  30'd    7171    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7172    : data = 32'h    014898B3    ;    //    sll x17 x17 x20      ====        sll a7, a7, s4
                                                  30'd    7173    : data = 32'h    B16D0493    ;    //    addi x9 x26 -1258      ====        addi s1, s10, -1258
                                                  30'd    7174    : data = 32'h    35C63DB7    ;    //    lui x27 220259      ====        lui s11, 220259
                                                  30'd    7175    : data = 32'h    714BA993    ;    //    slti x19 x23 1812      ====        slti s3, s7, 1812
                                                  30'd    7176    : data = 32'h    21F1A713    ;    //    slti x14 x3 543      ====        slti a4, gp, 543
                                                  30'd    7177    : data = 32'h    78C61897    ;    //    auipc x17 494689      ====        auipc a7, 494689
                                                  30'd    7178    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7179    : data = 32'h    40FDD133    ;    //    sra x2 x27 x15      ====        sra sp, s11, a5
                                                  30'd    7180    : data = 32'h    40445713    ;    //    srai x14 x8 4      ====        srai a4, s0, 4
                                                  30'd    7181    : data = 32'h    00ED98B3    ;    //    sll x17 x27 x14      ====        sll a7, s11, a4
                                                  30'd    7182    : data = 32'h    00A623B3    ;    //    slt x7 x12 x10      ====        slt t2, a2, a0
                                                  30'd    7183    : data = 32'h    007CE033    ;    //    or x0 x25 x7      ====        or zero, s9, t2
                                                  30'd    7184    : data = 32'h    6D432713    ;    //    slti x14 x6 1748      ====        slti a4, t1, 1748
                                                  30'd    7185    : data = 32'h    01DFE093    ;    //    ori x1 x31 29      ====        ori ra, t6, 29
                                                  30'd    7186    : data = 32'h    0194E6B3    ;    //    or x13 x9 x25      ====        or a3, s1, s9
                                                  30'd    7187    : data = 32'h    013CA333    ;    //    slt x6 x25 x19      ====        slt t1, s9, s3
                                                  30'd    7188    : data = 32'h    3A1C6F93    ;    //    ori x31 x24 929      ====        ori t6, s8, 929
                                                  30'd    7189    : data = 32'h    11122613    ;    //    slti x12 x4 273      ====        slti a2, tp, 273
                                                  30'd    7190    : data = 32'h    38AA2493    ;    //    slti x9 x20 906      ====        slti s1, s4, 906
                                                  30'd    7191    : data = 32'h    57596E13    ;    //    ori x28 x18 1397      ====        ori t3, s2, 1397
                                                  30'd    7192    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7193    : data = 32'h    97B00E93    ;    //    addi x29 x0 -1669      ====        addi t4, zero, -1669
                                                  30'd    7194    : data = 32'h    41DAD0B3    ;    //    sra x1 x21 x29      ====        sra ra, s5, t4
                                                  30'd    7195    : data = 32'h    418806B3    ;    //    sub x13 x16 x24      ====        sub a3, a6, s8
                                                  30'd    7196    : data = 32'h    77C67B93    ;    //    andi x23 x12 1916      ====        andi s7, a2, 1916
                                                  30'd    7197    : data = 32'h    01BD79B3    ;    //    and x19 x26 x27      ====        and s3, s10, s11
                                                  30'd    7198    : data = 32'h    165AF013    ;    //    andi x0 x21 357      ====        andi zero, s5, 357
                                                  30'd    7199    : data = 32'h    00928BB3    ;    //    add x23 x5 x9      ====        add s7, t0, s1
                                                  30'd    7200    : data = 32'h    58F57893    ;    //    andi x17 x10 1423      ====        andi a7, a0, 1423
                                                  30'd    7201    : data = 32'h    A4B32C13    ;    //    slti x24 x6 -1461      ====        slti s8, t1, -1461
                                                  30'd    7202    : data = 32'h    0E9791B7    ;    //    lui x3 59769      ====        lui gp, 59769
                                                  30'd    7203    : data = 32'h    56CEEE93    ;    //    ori x29 x29 1388      ====        ori t4, t4, 1388
                                                  30'd    7204    : data = 32'h    306F7B93    ;    //    andi x23 x30 774      ====        andi s7, t5, 774
                                                  30'd    7205    : data = 32'h    18642B37    ;    //    lui x22 99906      ====        lui s6, 99906
                                                  30'd    7206    : data = 32'h    013DDA13    ;    //    srli x20 x27 19      ====        srli s4, s11, 19
                                                  30'd    7207    : data = 32'h    D6FBF493    ;    //    andi x9 x23 -657      ====        andi s1, s7, -657
                                                  30'd    7208    : data = 32'h    011D26B3    ;    //    slt x13 x26 x17      ====        slt a3, s10, a7
                                                  30'd    7209    : data = 32'h    017531B3    ;    //    sltu x3 x10 x23      ====        sltu gp, a0, s7
                                                  30'd    7210    : data = 32'h    00A03D33    ;    //    sltu x26 x0 x10      ====        sltu s10, zero, a0
                                                  30'd    7211    : data = 32'h    CC792F93    ;    //    slti x31 x18 -825      ====        slti t6, s2, -825
                                                  30'd    7212    : data = 32'h    01E85B13    ;    //    srli x22 x16 30      ====        srli s6, a6, 30
                                                  30'd    7213    : data = 32'h    0113B4B3    ;    //    sltu x9 x7 x17      ====        sltu s1, t2, a7
                                                  30'd    7214    : data = 32'h    95CDB013    ;    //    sltiu x0 x27 -1700      ====        sltiu zero, s11, -1700
                                                  30'd    7215    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7216    : data = 32'h    03834FB7    ;    //    lui x31 14388      ====        lui t6, 14388
                                                  30'd    7217    : data = 32'h    22C77B97    ;    //    auipc x23 142455      ====        auipc s7, 142455
                                                  30'd    7218    : data = 32'h    DCC82D17    ;    //    auipc x26 904322      ====        auipc s10, 904322
                                                  30'd    7219    : data = 32'h    00FAD393    ;    //    srli x7 x21 15      ====        srli t2, s5, 15
                                                  30'd    7220    : data = 32'h    0040D693    ;    //    srli x13 x1 4      ====        srli a3, ra, 4
                                                  30'd    7221    : data = 32'h    01F49933    ;    //    sll x18 x9 x31      ====        sll s2, s1, t6
                                                  30'd    7222    : data = 32'h    5B559337    ;    //    lui x6 374105      ====        lui t1, 374105
                                                  30'd    7223    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7224    : data = 32'h    0016D793    ;    //    srli x15 x13 1      ====        srli a5, a3, 1
                                                  30'd    7225    : data = 32'h    2116AD13    ;    //    slti x26 x13 529      ====        slti s10, a3, 529
                                                  30'd    7226    : data = 32'h    C53964B7    ;    //    lui x9 807830      ====        lui s1, 807830
                                                  30'd    7227    : data = 32'h    9E21C093    ;    //    xori x1 x3 -1566      ====        xori ra, gp, -1566
                                                  30'd    7228    : data = 32'h    805BCA13    ;    //    xori x20 x23 -2043      ====        xori s4, s7, -2043
                                                  30'd    7229    : data = 32'h    4062D193    ;    //    srai x3 x5 6      ====        srai gp, t0, 6
                                                  30'd    7230    : data = 32'h    015F90B3    ;    //    sll x1 x31 x21      ====        sll ra, t6, s5
                                                  30'd    7231    : data = 32'h    003257B3    ;    //    srl x15 x4 x3      ====        srl a5, tp, gp
                                                  30'd    7232    : data = 32'h    002C41B3    ;    //    xor x3 x24 x2      ====        xor gp, s8, sp
                                                  30'd    7233    : data = 32'h    8CA06A13    ;    //    ori x20 x0 -1846      ====        ori s4, zero, -1846
                                                  30'd    7234    : data = 32'h    000C71B3    ;    //    and x3 x24 x0      ====        and gp, s8, zero
                                                  30'd    7235    : data = 32'h    BD9F8B97    ;    //    auipc x23 776696      ====        auipc s7, 776696
                                                  30'd    7236    : data = 32'h    012B5933    ;    //    srl x18 x22 x18      ====        srl s2, s6, s2
                                                  30'd    7237    : data = 32'h    40EC57B3    ;    //    sra x15 x24 x14      ====        sra a5, s8, a4
                                                  30'd    7238    : data = 32'h    014D63B3    ;    //    or x7 x26 x20      ====        or t2, s10, s4
                                                  30'd    7239    : data = 32'h    00299E33    ;    //    sll x28 x19 x2      ====        sll t3, s3, sp
                                                  30'd    7240    : data = 32'h    DCB1B937    ;    //    lui x18 903963      ====        lui s2, 903963
                                                  30'd    7241    : data = 32'h    E9F00D93    ;    //    addi x27 x0 -353      ====        addi s11, zero, -353
                                                  30'd    7242    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7243    : data = 32'h    00B39B33    ;    //    sll x22 x7 x11      ====        sll s6, t2, a1
                                                  30'd    7244    : data = 32'h    01C66833    ;    //    or x16 x12 x28      ====        or a6, a2, t3
                                                  30'd    7245    : data = 32'h    A3307D17    ;    //    auipc x26 668423      ====        auipc s10, 668423
                                                  30'd    7246    : data = 32'h    29A80913    ;    //    addi x18 x16 666      ====        addi s2, a6, 666
                                                  30'd    7247    : data = 32'h    2285CC93    ;    //    xori x25 x11 552      ====        xori s9, a1, 552
                                                  30'd    7248    : data = 32'h    A100FB13    ;    //    andi x22 x1 -1520      ====        andi s6, ra, -1520
                                                  30'd    7249    : data = 32'h    4951E313    ;    //    ori x6 x3 1173      ====        ori t1, gp, 1173
                                                  30'd    7250    : data = 32'h    9EE53337    ;    //    lui x6 650835      ====        lui t1, 650835
                                                  30'd    7251    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7252    : data = 32'h    006585B3    ;    //    add x11 x11 x6      ====        add a1, a1, t1
                                                  30'd    7253    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7254    : data = 32'h    14536713    ;    //    ori x14 x6 325      ====        ori a4, t1, 325
                                                  30'd    7255    : data = 32'h    CFB28E13    ;    //    addi x28 x5 -773      ====        addi t3, t0, -773
                                                  30'd    7256    : data = 32'h    002552B3    ;    //    srl x5 x10 x2      ====        srl t0, a0, sp
                                                  30'd    7257    : data = 32'h    402F06B3    ;    //    sub x13 x30 x2      ====        sub a3, t5, sp
                                                  30'd    7258    : data = 32'h    00FC30B3    ;    //    sltu x1 x24 x15      ====        sltu ra, s8, a5
                                                  30'd    7259    : data = 32'h    001F4B33    ;    //    xor x22 x30 x1      ====        xor s6, t5, ra
                                                  30'd    7260    : data = 32'h    00D3A333    ;    //    slt x6 x7 x13      ====        slt t1, t2, a3
                                                  30'd    7261    : data = 32'h    41D008B3    ;    //    sub x17 x0 x29      ====        sub a7, zero, t4
                                                  30'd    7262    : data = 32'h    40295F93    ;    //    srai x31 x18 2      ====        srai t6, s2, 2
                                                  30'd    7263    : data = 32'h    6EF87C13    ;    //    andi x24 x16 1775      ====        andi s8, a6, 1775
                                                  30'd    7264    : data = 32'h    0D8E6E97    ;    //    auipc x29 55526      ====        auipc t4, 55526
                                                  30'd    7265    : data = 32'h    6FE93613    ;    //    sltiu x12 x18 1790      ====        sltiu a2, s2, 1790
                                                  30'd    7266    : data = 32'h    400F89B3    ;    //    sub x19 x31 x0      ====        sub s3, t6, zero
                                                  30'd    7267    : data = 32'h    01B1FEB3    ;    //    and x29 x3 x27      ====        and t4, gp, s11
                                                  30'd    7268    : data = 32'h    00A876B3    ;    //    and x13 x16 x10      ====        and a3, a6, a0
                                                  30'd    7269    : data = 32'h    01B1D393    ;    //    srli x7 x3 27      ====        srli t2, gp, 27
                                                  30'd    7270    : data = 32'h    01A0D833    ;    //    srl x16 x1 x26      ====        srl a6, ra, s10
                                                  30'd    7271    : data = 32'h    40608093    ;    //    addi x1 x1 1030      ====        addi ra, ra, 1030
                                                  30'd    7272    : data = 32'h    009C21B3    ;    //    slt x3 x24 x9      ====        slt gp, s8, s1
                                                  30'd    7273    : data = 32'h    DD2F8293    ;    //    addi x5 x31 -558      ====        addi t0, t6, -558
                                                  30'd    7274    : data = 32'h    3FFEAA13    ;    //    slti x20 x29 1023      ====        slti s4, t4, 1023
                                                  30'd    7275    : data = 32'h    40D853B3    ;    //    sra x7 x16 x13      ====        sra t2, a6, a3
                                                  30'd    7276    : data = 32'h    01CF2B33    ;    //    slt x22 x30 x28      ====        slt s6, t5, t3
                                                  30'd    7277    : data = 32'h    4E0FE593    ;    //    ori x11 x31 1248      ====        ori a1, t6, 1248
                                                  30'd    7278    : data = 32'h    E9513117    ;    //    auipc x2 955667      ====        auipc sp, 955667
                                                  30'd    7279    : data = 32'h    00042A33    ;    //    slt x20 x8 x0      ====        slt s4, s0, zero
                                                  30'd    7280    : data = 32'h    47ABA413    ;    //    slti x8 x23 1146      ====        slti s0, s7, 1146
                                                  30'd    7281    : data = 32'h    40B35413    ;    //    srai x8 x6 11      ====        srai s0, t1, 11
                                                  30'd    7282    : data = 32'h    00F0F5B3    ;    //    and x11 x1 x15      ====        and a1, ra, a5
                                                  30'd    7283    : data = 32'h    00F530B3    ;    //    sltu x1 x10 x15      ====        sltu ra, a0, a5
                                                  30'd    7284    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7285    : data = 32'h    DBB8C693    ;    //    xori x13 x17 -581      ====        xori a3, a7, -581
                                                  30'd    7286    : data = 32'h    9C47AF93    ;    //    slti x31 x15 -1596      ====        slti t6, a5, -1596
                                                  30'd    7287    : data = 32'h    01654733    ;    //    xor x14 x10 x22      ====        xor a4, a0, s6
                                                  30'd    7288    : data = 32'h    24C92893    ;    //    slti x17 x18 588      ====        slti a7, s2, 588
                                                  30'd    7289    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7290    : data = 32'h    41A759B3    ;    //    sra x19 x14 x26      ====        sra s3, a4, s10
                                                  30'd    7291    : data = 32'h    014122B3    ;    //    slt x5 x2 x20      ====        slt t0, sp, s4
                                                  30'd    7292    : data = 32'h    44684113    ;    //    xori x2 x16 1094      ====        xori sp, a6, 1094
                                                  30'd    7293    : data = 32'h    01CE59B3    ;    //    srl x19 x28 x28      ====        srl s3, t3, t3
                                                  30'd    7294    : data = 32'h    00C867B3    ;    //    or x15 x16 x12      ====        or a5, a6, a2
                                                  30'd    7295    : data = 32'h    00F087B3    ;    //    add x15 x1 x15      ====        add a5, ra, a5
                                                  30'd    7296    : data = 32'h    00FA4D33    ;    //    xor x26 x20 x15      ====        xor s10, s4, a5
                                                  30'd    7297    : data = 32'h    008D5193    ;    //    srli x3 x26 8      ====        srli gp, s10, 8
                                                  30'd    7298    : data = 32'h    03753B13    ;    //    sltiu x22 x10 55      ====        sltiu s6, a0, 55
                                                  30'd    7299    : data = 32'h    008B7CB3    ;    //    and x25 x22 x8      ====        and s9, s6, s0
                                                  30'd    7300    : data = 32'h    41BD0EB3    ;    //    sub x29 x26 x27      ====        sub t4, s10, s11
                                                  30'd    7301    : data = 32'h    40EC89B3    ;    //    sub x19 x25 x14      ====        sub s3, s9, a4
                                                  30'd    7302    : data = 32'h    0069D313    ;    //    srli x6 x19 6      ====        srli t1, s3, 6
                                                  30'd    7303    : data = 32'h    0044E033    ;    //    or x0 x9 x4      ====        or zero, s1, tp
                                                  30'd    7304    : data = 32'h    40E75E93    ;    //    srai x29 x14 14      ====        srai t4, a4, 14
                                                  30'd    7305    : data = 32'h    00949FB3    ;    //    sll x31 x9 x9      ====        sll t6, s1, s1
                                                  30'd    7306    : data = 32'h    01D78833    ;    //    add x16 x15 x29      ====        add a6, a5, t4
                                                  30'd    7307    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7308    : data = 32'h    00ACD813    ;    //    srli x16 x25 10      ====        srli a6, s9, 10
                                                  30'd    7309    : data = 32'h    3B1A7493    ;    //    andi x9 x20 945      ====        andi s1, s4, 945
                                                  30'd    7310    : data = 32'h    007A6633    ;    //    or x12 x20 x7      ====        or a2, s4, t2
                                                  30'd    7311    : data = 32'h    411C5A33    ;    //    sra x20 x24 x17      ====        sra s4, s8, a7
                                                  30'd    7312    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7313    : data = 32'h    86199497    ;    //    auipc x9 549273      ====        auipc s1, 549273
                                                  30'd    7314    : data = 32'h    01348033    ;    //    add x0 x9 x19      ====        add zero, s1, s3
                                                  30'd    7315    : data = 32'h    00FA1D93    ;    //    slli x27 x20 15      ====        slli s11, s4, 15
                                                  30'd    7316    : data = 32'h    00665993    ;    //    srli x19 x12 6      ====        srli s3, a2, 6
                                                  30'd    7317    : data = 32'h    0149CA33    ;    //    xor x20 x19 x20      ====        xor s4, s3, s4
                                                  30'd    7318    : data = 32'h    563EE313    ;    //    ori x6 x29 1379      ====        ori t1, t4, 1379
                                                  30'd    7319    : data = 32'h    00BED593    ;    //    srli x11 x29 11      ====        srli a1, t4, 11
                                                  30'd    7320    : data = 32'h    01B6D7B3    ;    //    srl x15 x13 x27      ====        srl a5, a3, s11
                                                  30'd    7321    : data = 32'h    64EE0913    ;    //    addi x18 x28 1614      ====        addi s2, t3, 1614
                                                  30'd    7322    : data = 32'h    01CAF333    ;    //    and x6 x21 x28      ====        and t1, s5, t3
                                                  30'd    7323    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7324    : data = 32'h    A0812613    ;    //    slti x12 x2 -1528      ====        slti a2, sp, -1528
                                                  30'd    7325    : data = 32'h    01305BB3    ;    //    srl x23 x0 x19      ====        srl s7, zero, s3
                                                  30'd    7326    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7327    : data = 32'h    01A4C433    ;    //    xor x8 x9 x26      ====        xor s0, s1, s10
                                                  30'd    7328    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7329    : data = 32'h    41B15AB3    ;    //    sra x21 x2 x27      ====        sra s5, sp, s11
                                                  30'd    7330    : data = 32'h    00BA5933    ;    //    srl x18 x20 x11      ====        srl s2, s4, a1
                                                  30'd    7331    : data = 32'h    005ED313    ;    //    srli x6 x29 5      ====        srli t1, t4, 5
                                                  30'd    7332    : data = 32'h    91DD0B97    ;    //    auipc x23 597456      ====        auipc s7, 597456
                                                  30'd    7333    : data = 32'h    17B38397    ;    //    auipc x7 97080      ====        auipc t2, 97080
                                                  30'd    7334    : data = 32'h    823DC193    ;    //    xori x3 x27 -2013      ====        xori gp, s11, -2013
                                                  30'd    7335    : data = 32'h    06126493    ;    //    ori x9 x4 97      ====        ori s1, tp, 97
                                                  30'd    7336    : data = 32'h    40C901B3    ;    //    sub x3 x18 x12      ====        sub gp, s2, a2
                                                  30'd    7337    : data = 32'h    00B2ACB3    ;    //    slt x25 x5 x11      ====        slt s9, t0, a1
                                                  30'd    7338    : data = 32'h    72AA2D13    ;    //    slti x26 x20 1834      ====        slti s10, s4, 1834
                                                  30'd    7339    : data = 32'h    013CC5B3    ;    //    xor x11 x25 x19      ====        xor a1, s9, s3
                                                  30'd    7340    : data = 32'h    01792DB3    ;    //    slt x27 x18 x23      ====        slt s11, s2, s7
                                                  30'd    7341    : data = 32'h    013D6133    ;    //    or x2 x26 x19      ====        or sp, s10, s3
                                                  30'd    7342    : data = 32'h    01F5A433    ;    //    slt x8 x11 x31      ====        slt s0, a1, t6
                                                  30'd    7343    : data = 32'h    007E6D33    ;    //    or x26 x28 x7      ====        or s10, t3, t2
                                                  30'd    7344    : data = 32'h    40F95393    ;    //    srai x7 x18 15      ====        srai t2, s2, 15
                                                  30'd    7345    : data = 32'h    E130C113    ;    //    xori x2 x1 -493      ====        xori sp, ra, -493
                                                  30'd    7346    : data = 32'h    412F52B3    ;    //    sra x5 x30 x18      ====        sra t0, t5, s2
                                                  30'd    7347    : data = 32'h    01569B13    ;    //    slli x22 x13 21      ====        slli s6, a3, 21
                                                  30'd    7348    : data = 32'h    0038A3B3    ;    //    slt x7 x17 x3      ====        slt t2, a7, gp
                                                  30'd    7349    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7350    : data = 32'h    40A8E637    ;    //    lui x12 264846      ====        lui a2, 264846
                                                  30'd    7351    : data = 32'h    011597B3    ;    //    sll x15 x11 x17      ====        sll a5, a1, a7
                                                  30'd    7352    : data = 32'h    006564B3    ;    //    or x9 x10 x6      ====        or s1, a0, t1
                                                  30'd    7353    : data = 32'h    DA742113    ;    //    slti x2 x8 -601      ====        slti sp, s0, -601
                                                  30'd    7354    : data = 32'h    F3693F97    ;    //    auipc x31 997011      ====        auipc t6, 997011
                                                  30'd    7355    : data = 32'h    00B1D033    ;    //    srl x0 x3 x11      ====        srl zero, gp, a1
                                                  30'd    7356    : data = 32'h    2654F693    ;    //    andi x13 x9 613      ====        andi a3, s1, 613
                                                  30'd    7357    : data = 32'h    002B64B3    ;    //    or x9 x22 x2      ====        or s1, s6, sp
                                                  30'd    7358    : data = 32'h    002FABB3    ;    //    slt x23 x31 x2      ====        slt s7, t6, sp
                                                  30'd    7359    : data = 32'h    4056D933    ;    //    sra x18 x13 x5      ====        sra s2, a3, t0
                                                  30'd    7360    : data = 32'h    41070133    ;    //    sub x2 x14 x16      ====        sub sp, a4, a6
                                                  30'd    7361    : data = 32'h    35582137    ;    //    lui x2 218498      ====        lui sp, 218498
                                                  30'd    7362    : data = 32'h    8F962713    ;    //    slti x14 x12 -1799      ====        slti a4, a2, -1799
                                                  30'd    7363    : data = 32'h    010FDBB3    ;    //    srl x23 x31 x16      ====        srl s7, t6, a6
                                                  30'd    7364    : data = 32'h    00E584B3    ;    //    add x9 x11 x14      ====        add s1, a1, a4
                                                  30'd    7365    : data = 32'h    97200997    ;    //    auipc x19 619008      ====        auipc s3, 619008
                                                  30'd    7366    : data = 32'h    EAB07713    ;    //    andi x14 x0 -341      ====        andi a4, zero, -341
                                                  30'd    7367    : data = 32'h    40210133    ;    //    sub x2 x2 x2      ====        sub sp, sp, sp
                                                  30'd    7368    : data = 32'h    94D4A713    ;    //    slti x14 x9 -1715      ====        slti a4, s1, -1715
                                                  30'd    7369    : data = 32'h    3BEA8D13    ;    //    addi x26 x21 958      ====        addi s10, s5, 958
                                                  30'd    7370    : data = 32'h    00B70333    ;    //    add x6 x14 x11      ====        add t1, a4, a1
                                                  30'd    7371    : data = 32'h    00342833    ;    //    slt x16 x8 x3      ====        slt a6, s0, gp
                                                  30'd    7372    : data = 32'h    011B1A13    ;    //    slli x20 x22 17      ====        slli s4, s6, 17
                                                  30'd    7373    : data = 32'h    0011E8B3    ;    //    or x17 x3 x1      ====        or a7, gp, ra
                                                  30'd    7374    : data = 32'h    7ECE9437    ;    //    lui x8 519401      ====        lui s0, 519401
                                                  30'd    7375    : data = 32'h    E2C0CD97    ;    //    auipc x27 928780      ====        auipc s11, 928780
                                                  30'd    7376    : data = 32'h    018EBAB3    ;    //    sltu x21 x29 x24      ====        sltu s5, t4, s8
                                                  30'd    7377    : data = 32'h    D204FA13    ;    //    andi x20 x9 -736      ====        andi s4, s1, -736
                                                  30'd    7378    : data = 32'h    70087993    ;    //    andi x19 x16 1792      ====        andi s3, a6, 1792
                                                  30'd    7379    : data = 32'h    405E5033    ;    //    sra x0 x28 x5      ====        sra zero, t3, t0
                                                  30'd    7380    : data = 32'h    01DFB833    ;    //    sltu x16 x31 x29      ====        sltu a6, t6, t4
                                                  30'd    7381    : data = 32'h    41590DB3    ;    //    sub x27 x18 x21      ====        sub s11, s2, s5
                                                  30'd    7382    : data = 32'h    ABD03693    ;    //    sltiu x13 x0 -1347      ====        sltiu a3, zero, -1347
                                                  30'd    7383    : data = 32'h    01ADF6B3    ;    //    and x13 x27 x26      ====        and a3, s11, s10
                                                  30'd    7384    : data = 32'h    40385433    ;    //    sra x8 x16 x3      ====        sra s0, a6, gp
                                                  30'd    7385    : data = 32'h    EC28AB13    ;    //    slti x22 x17 -318      ====        slti s6, a7, -318
                                                  30'd    7386    : data = 32'h    A568CB93    ;    //    xori x23 x17 -1450      ====        xori s7, a7, -1450
                                                  30'd    7387    : data = 32'h    0115AC33    ;    //    slt x24 x11 x17      ====        slt s8, a1, a7
                                                  30'd    7388    : data = 32'h    41358FB3    ;    //    sub x31 x11 x19      ====        sub t6, a1, s3
                                                  30'd    7389    : data = 32'h    F941EE93    ;    //    ori x29 x3 -108      ====        ori t4, gp, -108
                                                  30'd    7390    : data = 32'h    0114F4B3    ;    //    and x9 x9 x17      ====        and s1, s1, a7
                                                  30'd    7391    : data = 32'h    AE3D4193    ;    //    xori x3 x26 -1309      ====        xori gp, s10, -1309
                                                  30'd    7392    : data = 32'h    01B422B3    ;    //    slt x5 x8 x27      ====        slt t0, s0, s11
                                                  30'd    7393    : data = 32'h    009849B3    ;    //    xor x19 x16 x9      ====        xor s3, a6, s1
                                                  30'd    7394    : data = 32'h    01C66933    ;    //    or x18 x12 x28      ====        or s2, a2, t3
                                                  30'd    7395    : data = 32'h    D17DE093    ;    //    ori x1 x27 -745      ====        ori ra, s11, -745
                                                  30'd    7396    : data = 32'h    01BC2CB3    ;    //    slt x25 x24 x27      ====        slt s9, s8, s11
                                                  30'd    7397    : data = 32'h    01465DB3    ;    //    srl x27 x12 x20      ====        srl s11, a2, s4
                                                  30'd    7398    : data = 32'h    00A628B3    ;    //    slt x17 x12 x10      ====        slt a7, a2, a0
                                                  30'd    7399    : data = 32'h    011A1893    ;    //    slli x17 x20 17      ====        slli a7, s4, 17
                                                  30'd    7400    : data = 32'h    404E0B33    ;    //    sub x22 x28 x4      ====        sub s6, t3, tp
                                                  30'd    7401    : data = 32'h    6503D837    ;    //    lui x16 413757      ====        lui a6, 413757
                                                  30'd    7402    : data = 32'h    7A17C613    ;    //    xori x12 x15 1953      ====        xori a2, a5, 1953
                                                  30'd    7403    : data = 32'h    D7B37A93    ;    //    andi x21 x6 -645      ====        andi s5, t1, -645
                                                  30'd    7404    : data = 32'h    E48741B7    ;    //    lui x3 936052      ====        lui gp, 936052
                                                  30'd    7405    : data = 32'h    0048A5B3    ;    //    slt x11 x17 x4      ====        slt a1, a7, tp
                                                  30'd    7406    : data = 32'h    BE9B8B93    ;    //    addi x23 x23 -1047      ====        addi s7, s7, -1047
                                                  30'd    7407    : data = 32'h    01928D33    ;    //    add x26 x5 x25      ====        add s10, t0, s9
                                                  30'd    7408    : data = 32'h    40B65613    ;    //    srai x12 x12 11      ====        srai a2, a2, 11
                                                  30'd    7409    : data = 32'h    E27DA717    ;    //    auipc x14 927706      ====        auipc a4, 927706
                                                  30'd    7410    : data = 32'h    D50B4693    ;    //    xori x13 x22 -688      ====        xori a3, s6, -688
                                                  30'd    7411    : data = 32'h    00BA70B3    ;    //    and x1 x20 x11      ====        and ra, s4, a1
                                                  30'd    7412    : data = 32'h    01A95633    ;    //    srl x12 x18 x26      ====        srl a2, s2, s10
                                                  30'd    7413    : data = 32'h    00CFDA93    ;    //    srli x21 x31 12      ====        srli s5, t6, 12
                                                  30'd    7414    : data = 32'h    011F1B33    ;    //    sll x22 x30 x17      ====        sll s6, t5, a7
                                                  30'd    7415    : data = 32'h    00753833    ;    //    sltu x16 x10 x7      ====        sltu a6, a0, t2
                                                  30'd    7416    : data = 32'h    01157033    ;    //    and x0 x10 x17      ====        and zero, a0, a7
                                                  30'd    7417    : data = 32'h    419A80B3    ;    //    sub x1 x21 x25      ====        sub ra, s5, s9
                                                  30'd    7418    : data = 32'h    76DEB013    ;    //    sltiu x0 x29 1901      ====        sltiu zero, t4, 1901
                                                  30'd    7419    : data = 32'h    012219B3    ;    //    sll x19 x4 x18      ====        sll s3, tp, s2
                                                  30'd    7420    : data = 32'h    B870D017    ;    //    auipc x0 755469      ====        auipc zero, 755469
                                                  30'd    7421    : data = 32'h    003A5B13    ;    //    srli x22 x20 3      ====        srli s6, s4, 3
                                                  30'd    7422    : data = 32'h    01769393    ;    //    slli x7 x13 23      ====        slli t2, a3, 23
                                                  30'd    7423    : data = 32'h    A1E6C993    ;    //    xori x19 x13 -1506      ====        xori s3, a3, -1506
                                                  30'd    7424    : data = 32'h    00A199B3    ;    //    sll x19 x3 x10      ====        sll s3, gp, a0
                                                  30'd    7425    : data = 32'h    FC9EA993    ;    //    slti x19 x29 -55      ====        slti s3, t4, -55
                                                  30'd    7426    : data = 32'h    007B56B3    ;    //    srl x13 x22 x7      ====        srl a3, s6, t2
                                                  30'd    7427    : data = 32'h    5CE67613    ;    //    andi x12 x12 1486      ====        andi a2, a2, 1486
                                                  30'd    7428    : data = 32'h    01499413    ;    //    slli x8 x19 20      ====        slli s0, s3, 20
                                                  30'd    7429    : data = 32'h    000C4AB3    ;    //    xor x21 x24 x0      ====        xor s5, s8, zero
                                                  30'd    7430    : data = 32'h    AE927E13    ;    //    andi x28 x4 -1303      ====        andi t3, tp, -1303
                                                  30'd    7431    : data = 32'h    0132AEB3    ;    //    slt x29 x5 x19      ====        slt t4, t0, s3
                                                  30'd    7432    : data = 32'h    00526433    ;    //    or x8 x4 x5      ====        or s0, tp, t0
                                                  30'd    7433    : data = 32'h    D1007993    ;    //    andi x19 x0 -752      ====        andi s3, zero, -752
                                                  30'd    7434    : data = 32'h    40978CB3    ;    //    sub x25 x15 x9      ====        sub s9, a5, s1
                                                  30'd    7435    : data = 32'h    B5E77013    ;    //    andi x0 x14 -1186      ====        andi zero, a4, -1186
                                                  30'd    7436    : data = 32'h    5290CA97    ;    //    auipc x21 338188      ====        auipc s5, 338188
                                                  30'd    7437    : data = 32'h    01859113    ;    //    slli x2 x11 24      ====        slli sp, a1, 24
                                                  30'd    7438    : data = 32'h    016536B3    ;    //    sltu x13 x10 x22      ====        sltu a3, a0, s6
                                                  30'd    7439    : data = 32'h    010B94B3    ;    //    sll x9 x23 x16      ====        sll s1, s7, a6
                                                  30'd    7440    : data = 32'h    31078413    ;    //    addi x8 x15 784      ====        addi s0, a5, 784
                                                  30'd    7441    : data = 32'h    010833B3    ;    //    sltu x7 x16 x16      ====        sltu t2, a6, a6
                                                  30'd    7442    : data = 32'h    4120D4B3    ;    //    sra x9 x1 x18      ====        sra s1, ra, s2
                                                  30'd    7443    : data = 32'h    0094CA33    ;    //    xor x20 x9 x9      ====        xor s4, s1, s1
                                                  30'd    7444    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7445    : data = 32'h    0024C633    ;    //    xor x12 x9 x2      ====        xor a2, s1, sp
                                                  30'd    7446    : data = 32'h    9ABB4897    ;    //    auipc x17 633780      ====        auipc a7, 633780
                                                  30'd    7447    : data = 32'h    01FA41B3    ;    //    xor x3 x20 x31      ====        xor gp, s4, t6
                                                  30'd    7448    : data = 32'h    005F6DB3    ;    //    or x27 x30 x5      ====        or s11, t5, t0
                                                  30'd    7449    : data = 32'h    40FE5BB3    ;    //    sra x23 x28 x15      ====        sra s7, t3, a5
                                                  30'd    7450    : data = 32'h    9838B413    ;    //    sltiu x8 x17 -1661      ====        sltiu s0, a7, -1661
                                                  30'd    7451    : data = 32'h    7B1F7013    ;    //    andi x0 x30 1969      ====        andi zero, t5, 1969
                                                  30'd    7452    : data = 32'h    0096E5B3    ;    //    or x11 x13 x9      ====        or a1, a3, s1
                                                  30'd    7453    : data = 32'h    0051B633    ;    //    sltu x12 x3 x5      ====        sltu a2, gp, t0
                                                  30'd    7454    : data = 32'h    332A7393    ;    //    andi x7 x20 818      ====        andi t2, s4, 818
                                                  30'd    7455    : data = 32'h    01CEBD33    ;    //    sltu x26 x29 x28      ====        sltu s10, t4, t3
                                                  30'd    7456    : data = 32'h    00D712B3    ;    //    sll x5 x14 x13      ====        sll t0, a4, a3
                                                  30'd    7457    : data = 32'h    E34C7E93    ;    //    andi x29 x24 -460      ====        andi t4, s8, -460
                                                  30'd    7458    : data = 32'h    010C1D93    ;    //    slli x27 x24 16      ====        slli s11, s8, 16
                                                  30'd    7459    : data = 32'h    01D68333    ;    //    add x6 x13 x29      ====        add t1, a3, t4
                                                  30'd    7460    : data = 32'h    00921A13    ;    //    slli x20 x4 9      ====        slli s4, tp, 9
                                                  30'd    7461    : data = 32'h    41D082B3    ;    //    sub x5 x1 x29      ====        sub t0, ra, t4
                                                  30'd    7462    : data = 32'h    C730AA13    ;    //    slti x20 x1 -909      ====        slti s4, ra, -909
                                                  30'd    7463    : data = 32'h    019B5413    ;    //    srli x8 x22 25      ====        srli s0, s6, 25
                                                  30'd    7464    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7465    : data = 32'h    F48BA913    ;    //    slti x18 x23 -184      ====        slti s2, s7, -184
                                                  30'd    7466    : data = 32'h    2A816797    ;    //    auipc x15 174102      ====        auipc a5, 174102
                                                  30'd    7467    : data = 32'h    41BADFB3    ;    //    sra x31 x21 x27      ====        sra t6, s5, s11
                                                  30'd    7468    : data = 32'h    00BD9333    ;    //    sll x6 x27 x11      ====        sll t1, s11, a1
                                                  30'd    7469    : data = 32'h    3583FE97    ;    //    auipc x29 219199      ====        auipc t4, 219199
                                                  30'd    7470    : data = 32'h    015F33B3    ;    //    sltu x7 x30 x21      ====        sltu t2, t5, s5
                                                  30'd    7471    : data = 32'h    410CDA13    ;    //    srai x20 x25 16      ====        srai s4, s9, 16
                                                  30'd    7472    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7473    : data = 32'h    015C7D33    ;    //    and x26 x24 x21      ====        and s10, s8, s5
                                                  30'd    7474    : data = 32'h    41788833    ;    //    sub x16 x17 x23      ====        sub a6, a7, s7
                                                  30'd    7475    : data = 32'h    015DEE33    ;    //    or x28 x27 x21      ====        or t3, s11, s5
                                                  30'd    7476    : data = 32'h    01B334B3    ;    //    sltu x9 x6 x27      ====        sltu s1, t1, s11
                                                  30'd    7477    : data = 32'h    BF9ABD13    ;    //    sltiu x26 x21 -1031      ====        sltiu s10, s5, -1031
                                                  30'd    7478    : data = 32'h    EE15E313    ;    //    ori x6 x11 -287      ====        ori t1, a1, -287
                                                  30'd    7479    : data = 32'h    000F5A13    ;    //    srli x20 x30 0      ====        srli s4, t5, 0
                                                  30'd    7480    : data = 32'h    013C70B3    ;    //    and x1 x24 x19      ====        and ra, s8, s3
                                                  30'd    7481    : data = 32'h    005F67B3    ;    //    or x15 x30 x5      ====        or a5, t5, t0
                                                  30'd    7482    : data = 32'h    FEA13C93    ;    //    sltiu x25 x2 -22      ====        sltiu s9, sp, -22
                                                  30'd    7483    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7484    : data = 32'h    4FB9A813    ;    //    slti x16 x19 1275      ====        slti a6, s3, 1275
                                                  30'd    7485    : data = 32'h    40EB8D33    ;    //    sub x26 x23 x14      ====        sub s10, s7, a4
                                                  30'd    7486    : data = 32'h    009D9993    ;    //    slli x19 x27 9      ====        slli s3, s11, 9
                                                  30'd    7487    : data = 32'h    01C03033    ;    //    sltu x0 x0 x28      ====        sltu zero, zero, t3
                                                  30'd    7488    : data = 32'h    002F6633    ;    //    or x12 x30 x2      ====        or a2, t5, sp
                                                  30'd    7489    : data = 32'h    01E41713    ;    //    slli x14 x8 30      ====        slli a4, s0, 30
                                                  30'd    7490    : data = 32'h    CB38BF97    ;    //    auipc x31 832395      ====        auipc t6, 832395
                                                  30'd    7491    : data = 32'h    00D19713    ;    //    slli x14 x3 13      ====        slli a4, gp, 13
                                                  30'd    7492    : data = 32'h    004A5CB3    ;    //    srl x25 x20 x4      ====        srl s9, s4, tp
                                                  30'd    7493    : data = 32'h    40D2DBB3    ;    //    sra x23 x5 x13      ====        sra s7, t0, a3
                                                  30'd    7494    : data = 32'h    00301893    ;    //    slli x17 x0 3      ====        slli a7, zero, 3
                                                  30'd    7495    : data = 32'h    FC270D13    ;    //    addi x26 x14 -62      ====        addi s10, a4, -62
                                                  30'd    7496    : data = 32'h    EB46AA13    ;    //    slti x20 x13 -332      ====        slti s4, a3, -332
                                                  30'd    7497    : data = 32'h    41E1DBB3    ;    //    sra x23 x3 x30      ====        sra s7, gp, t5
                                                  30'd    7498    : data = 32'h    40ACD333    ;    //    sra x6 x25 x10      ====        sra t1, s9, a0
                                                  30'd    7499    : data = 32'h    66C22313    ;    //    slti x6 x4 1644      ====        slti t1, tp, 1644
                                                  30'd    7500    : data = 32'h    F5B18493    ;    //    addi x9 x3 -165      ====        addi s1, gp, -165
                                                  30'd    7501    : data = 32'h    AF30EA13    ;    //    ori x20 x1 -1293      ====        ori s4, ra, -1293
                                                  30'd    7502    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7503    : data = 32'h    01AAC833    ;    //    xor x16 x21 x26      ====        xor a6, s5, s10
                                                  30'd    7504    : data = 32'h    00622C33    ;    //    slt x24 x4 x6      ====        slt s8, tp, t1
                                                  30'd    7505    : data = 32'h    2EB26013    ;    //    ori x0 x4 747      ====        ori zero, tp, 747
                                                  30'd    7506    : data = 32'h    D887B3B7    ;    //    lui x7 886907      ====        lui t2, 886907
                                                  30'd    7507    : data = 32'h    B07E7693    ;    //    andi x13 x28 -1273      ====        andi a3, t3, -1273
                                                  30'd    7508    : data = 32'h    01B64EB3    ;    //    xor x29 x12 x27      ====        xor t4, a2, s11
                                                  30'd    7509    : data = 32'h    003A1993    ;    //    slli x19 x20 3      ====        slli s3, s4, 3
                                                  30'd    7510    : data = 32'h    34F9CB13    ;    //    xori x22 x19 847      ====        xori s6, s3, 847
                                                  30'd    7511    : data = 32'h    00FB8C33    ;    //    add x24 x23 x15      ====        add s8, s7, a5
                                                  30'd    7512    : data = 32'h    01462D33    ;    //    slt x26 x12 x20      ====        slt s10, a2, s4
                                                  30'd    7513    : data = 32'h    8E8ABC13    ;    //    sltiu x24 x21 -1816      ====        sltiu s8, s5, -1816
                                                  30'd    7514    : data = 32'h    00E95433    ;    //    srl x8 x18 x14      ====        srl s0, s2, a4
                                                  30'd    7515    : data = 32'h    0087D933    ;    //    srl x18 x15 x8      ====        srl s2, a5, s0
                                                  30'd    7516    : data = 32'h    40585C33    ;    //    sra x24 x16 x5      ====        sra s8, a6, t0
                                                  30'd    7517    : data = 32'h    16950393    ;    //    addi x7 x10 361      ====        addi t2, a0, 361
                                                  30'd    7518    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7519    : data = 32'h    00978EB3    ;    //    add x29 x15 x9      ====        add t4, a5, s1
                                                  30'd    7520    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7521    : data = 32'h    0FAD7D97    ;    //    auipc x27 64215      ====        auipc s11, 64215
                                                  30'd    7522    : data = 32'h    00FE71B3    ;    //    and x3 x28 x15      ====        and gp, t3, a5
                                                  30'd    7523    : data = 32'h    40475133    ;    //    sra x2 x14 x4      ====        sra sp, a4, tp
                                                  30'd    7524    : data = 32'h    00FEA133    ;    //    slt x2 x29 x15      ====        slt sp, t4, a5
                                                  30'd    7525    : data = 32'h    013AC8B3    ;    //    xor x17 x21 x19      ====        xor a7, s5, s3
                                                  30'd    7526    : data = 32'h    31EA4C93    ;    //    xori x25 x20 798      ====        xori s9, s4, 798
                                                  30'd    7527    : data = 32'h    0048BC33    ;    //    sltu x24 x17 x4      ====        sltu s8, a7, tp
                                                  30'd    7528    : data = 32'h    01CDD793    ;    //    srli x15 x27 28      ====        srli a5, s11, 28
                                                  30'd    7529    : data = 32'h    0150CBB3    ;    //    xor x23 x1 x21      ====        xor s7, ra, s5
                                                  30'd    7530    : data = 32'h    4105D933    ;    //    sra x18 x11 x16      ====        sra s2, a1, a6
                                                  30'd    7531    : data = 32'h    00738BB3    ;    //    add x23 x7 x7      ====        add s7, t2, t2
                                                  30'd    7532    : data = 32'h    40345033    ;    //    sra x0 x8 x3      ====        sra zero, s0, gp
                                                  30'd    7533    : data = 32'h    00E9DC13    ;    //    srli x24 x19 14      ====        srli s8, s3, 14
                                                  30'd    7534    : data = 32'h    35AFAC13    ;    //    slti x24 x31 858      ====        slti s8, t6, 858
                                                  30'd    7535    : data = 32'h    00D365B3    ;    //    or x11 x6 x13      ====        or a1, t1, a3
                                                  30'd    7536    : data = 32'h    5B92BA93    ;    //    sltiu x21 x5 1465      ====        sltiu s5, t0, 1465
                                                  30'd    7537    : data = 32'h    01D15613    ;    //    srli x12 x2 29      ====        srli a2, sp, 29
                                                  30'd    7538    : data = 32'h    348FD897    ;    //    auipc x17 215293      ====        auipc a7, 215293
                                                  30'd    7539    : data = 32'h    000436B3    ;    //    sltu x13 x8 x0      ====        sltu a3, s0, zero
                                                  30'd    7540    : data = 32'h    00C9CB33    ;    //    xor x22 x19 x12      ====        xor s6, s3, a2
                                                  30'd    7541    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7542    : data = 32'h    059BE713    ;    //    ori x14 x23 89      ====        ori a4, s7, 89
                                                  30'd    7543    : data = 32'h    40A95613    ;    //    srai x12 x18 10      ====        srai a2, s2, 10
                                                  30'd    7544    : data = 32'h    01808B33    ;    //    add x22 x1 x24      ====        add s6, ra, s8
                                                  30'd    7545    : data = 32'h    0050FCB3    ;    //    and x25 x1 x5      ====        and s9, ra, t0
                                                  30'd    7546    : data = 32'h    00BC1413    ;    //    slli x8 x24 11      ====        slli s0, s8, 11
                                                  30'd    7547    : data = 32'h    95C54993    ;    //    xori x19 x10 -1700      ====        xori s3, a0, -1700
                                                  30'd    7548    : data = 32'h    01A75A33    ;    //    srl x20 x14 x26      ====        srl s4, a4, s10
                                                  30'd    7549    : data = 32'h    01E22733    ;    //    slt x14 x4 x30      ====        slt a4, tp, t5
                                                  30'd    7550    : data = 32'h    0000F2B3    ;    //    and x5 x1 x0      ====        and t0, ra, zero
                                                  30'd    7551    : data = 32'h    E216AB93    ;    //    slti x23 x13 -479      ====        slti s7, a3, -479
                                                  30'd    7552    : data = 32'h    BC762D13    ;    //    slti x26 x12 -1081      ====        slti s10, a2, -1081
                                                  30'd    7553    : data = 32'h    69413493    ;    //    sltiu x9 x2 1684      ====        sltiu s1, sp, 1684
                                                  30'd    7554    : data = 32'h    541F0413    ;    //    addi x8 x30 1345      ====        addi s0, t5, 1345
                                                  30'd    7555    : data = 32'h    8585BC93    ;    //    sltiu x25 x11 -1960      ====        sltiu s9, a1, -1960
                                                  30'd    7556    : data = 32'h    8D1EC413    ;    //    xori x8 x29 -1839      ====        xori s0, t4, -1839
                                                  30'd    7557    : data = 32'h    01C609B3    ;    //    add x19 x12 x28      ====        add s3, a2, t3
                                                  30'd    7558    : data = 32'h    C4C58713    ;    //    addi x14 x11 -948      ====        addi a4, a1, -948
                                                  30'd    7559    : data = 32'h    01B63033    ;    //    sltu x0 x12 x27      ====        sltu zero, a2, s11
                                                  30'd    7560    : data = 32'h    6098BA13    ;    //    sltiu x20 x17 1545      ====        sltiu s4, a7, 1545
                                                  30'd    7561    : data = 32'h    00D61933    ;    //    sll x18 x12 x13      ====        sll s2, a2, a3
                                                  30'd    7562    : data = 32'h    408F5133    ;    //    sra x2 x30 x8      ====        sra sp, t5, s0
                                                  30'd    7563    : data = 32'h    40A15A33    ;    //    sra x20 x2 x10      ====        sra s4, sp, a0
                                                  30'd    7564    : data = 32'h    00660833    ;    //    add x16 x12 x6      ====        add a6, a2, t1
                                                  30'd    7565    : data = 32'h    47B90113    ;    //    addi x2 x18 1147      ====        addi sp, s2, 1147
                                                  30'd    7566    : data = 32'h    00DF8E33    ;    //    add x28 x31 x13      ====        add t3, t6, a3
                                                  30'd    7567    : data = 32'h    00D1FAB3    ;    //    and x21 x3 x13      ====        and s5, gp, a3
                                                  30'd    7568    : data = 32'h    9DB08693    ;    //    addi x13 x1 -1573      ====        addi a3, ra, -1573
                                                  30'd    7569    : data = 32'h    0B704F93    ;    //    xori x31 x0 183      ====        xori t6, zero, 183
                                                  30'd    7570    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7571    : data = 32'h    00F19EB3    ;    //    sll x29 x3 x15      ====        sll t4, gp, a5
                                                  30'd    7572    : data = 32'h    40D7D7B3    ;    //    sra x15 x15 x13      ====        sra a5, a5, a3
                                                  30'd    7573    : data = 32'h    011F6D33    ;    //    or x26 x30 x17      ====        or s10, t5, a7
                                                  30'd    7574    : data = 32'h    00A67C33    ;    //    and x24 x12 x10      ====        and s8, a2, a0
                                                  30'd    7575    : data = 32'h    23D3E713    ;    //    ori x14 x7 573      ====        ori a4, t2, 573
                                                  30'd    7576    : data = 32'h    01C27A33    ;    //    and x20 x4 x28      ====        and s4, tp, t3
                                                  30'd    7577    : data = 32'h    01C76433    ;    //    or x8 x14 x28      ====        or s0, a4, t3
                                                  30'd    7578    : data = 32'h    D8C0E593    ;    //    ori x11 x1 -628      ====        ori a1, ra, -628
                                                  30'd    7579    : data = 32'h    55242593    ;    //    slti x11 x8 1362      ====        slti a1, s0, 1362
                                                  30'd    7580    : data = 32'h    01AC0933    ;    //    add x18 x24 x26      ====        add s2, s8, s10
                                                  30'd    7581    : data = 32'h    00E0ECB3    ;    //    or x25 x1 x14      ====        or s9, ra, a4
                                                  30'd    7582    : data = 32'h    E2D2E593    ;    //    ori x11 x5 -467      ====        ori a1, t0, -467
                                                  30'd    7583    : data = 32'h    01AF1033    ;    //    sll x0 x30 x26      ====        sll zero, t5, s10
                                                  30'd    7584    : data = 32'h    01B09F93    ;    //    slli x31 x1 27      ====        slli t6, ra, 27
                                                  30'd    7585    : data = 32'h    462C6993    ;    //    ori x19 x24 1122      ====        ori s3, s8, 1122
                                                  30'd    7586    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7587    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7588    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7589    : data = 32'h    413ED193    ;    //    srai x3 x29 19      ====        srai gp, t4, 19
                                                  30'd    7590    : data = 32'h    403C5893    ;    //    srai x17 x24 3      ====        srai a7, s8, 3
                                                  30'd    7591    : data = 32'h    2881F793    ;    //    andi x15 x3 648      ====        andi a5, gp, 648
                                                  30'd    7592    : data = 32'h    401FD6B3    ;    //    sra x13 x31 x1      ====        sra a3, t6, ra
                                                  30'd    7593    : data = 32'h    99BA3113    ;    //    sltiu x2 x20 -1637      ====        sltiu sp, s4, -1637
                                                  30'd    7594    : data = 32'h    01ADDB93    ;    //    srli x23 x27 26      ====        srli s7, s11, 26
                                                  30'd    7595    : data = 32'h    A516B193    ;    //    sltiu x3 x13 -1455      ====        sltiu gp, a3, -1455
                                                  30'd    7596    : data = 32'h    0190DCB3    ;    //    srl x25 x1 x25      ====        srl s9, ra, s9
                                                  30'd    7597    : data = 32'h    2EBBAD13    ;    //    slti x26 x23 747      ====        slti s10, s7, 747
                                                  30'd    7598    : data = 32'h    D271B413    ;    //    sltiu x8 x3 -729      ====        sltiu s0, gp, -729
                                                  30'd    7599    : data = 32'h    001EBCB3    ;    //    sltu x25 x29 x1      ====        sltu s9, t4, ra
                                                  30'd    7600    : data = 32'h    1BFB8713    ;    //    addi x14 x23 447      ====        addi a4, s7, 447
                                                  30'd    7601    : data = 32'h    411BD813    ;    //    srai x16 x23 17      ====        srai a6, s7, 17
                                                  30'd    7602    : data = 32'h    05912817    ;    //    auipc x16 22802      ====        auipc a6, 22802
                                                  30'd    7603    : data = 32'h    000C0733    ;    //    add x14 x24 x0      ====        add a4, s8, zero
                                                  30'd    7604    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7605    : data = 32'h    00C11FB3    ;    //    sll x31 x2 x12      ====        sll t6, sp, a2
                                                  30'd    7606    : data = 32'h    C3AA3E13    ;    //    sltiu x28 x20 -966      ====        sltiu t3, s4, -966
                                                  30'd    7607    : data = 32'h    419F0FB3    ;    //    sub x31 x30 x25      ====        sub t6, t5, s9
                                                  30'd    7608    : data = 32'h    01A0AFB3    ;    //    slt x31 x1 x26      ====        slt t6, ra, s10
                                                  30'd    7609    : data = 32'h    EE180693    ;    //    addi x13 x16 -287      ====        addi a3, a6, -287
                                                  30'd    7610    : data = 32'h    52E33413    ;    //    sltiu x8 x6 1326      ====        sltiu s0, t1, 1326
                                                  30'd    7611    : data = 32'h    413C0033    ;    //    sub x0 x24 x19      ====        sub zero, s8, s3
                                                  30'd    7612    : data = 32'h    00F051B3    ;    //    srl x3 x0 x15      ====        srl gp, zero, a5
                                                  30'd    7613    : data = 32'h    005ADC13    ;    //    srli x24 x21 5      ====        srli s8, s5, 5
                                                  30'd    7614    : data = 32'h    41F1BC93    ;    //    sltiu x25 x3 1055      ====        sltiu s9, gp, 1055
                                                  30'd    7615    : data = 32'h    0013DEB3    ;    //    srl x29 x7 x1      ====        srl t4, t2, ra
                                                  30'd    7616    : data = 32'h    011CAEB3    ;    //    slt x29 x25 x17      ====        slt t4, s9, a7
                                                  30'd    7617    : data = 32'h    4130D933    ;    //    sra x18 x1 x19      ====        sra s2, ra, s3
                                                  30'd    7618    : data = 32'h    00AC90B3    ;    //    sll x1 x25 x10      ====        sll ra, s9, a0
                                                  30'd    7619    : data = 32'h    73F2C913    ;    //    xori x18 x5 1855      ====        xori s2, t0, 1855
                                                  30'd    7620    : data = 32'h    759C8293    ;    //    addi x5 x25 1881      ====        addi t0, s9, 1881
                                                  30'd    7621    : data = 32'h    EFB30993    ;    //    addi x19 x6 -261      ====        addi s3, t1, -261
                                                  30'd    7622    : data = 32'h    40585593    ;    //    srai x11 x16 5      ====        srai a1, a6, 5
                                                  30'd    7623    : data = 32'h    01FB0133    ;    //    add x2 x22 x31      ====        add sp, s6, t6
                                                  30'd    7624    : data = 32'h    009A05B3    ;    //    add x11 x20 x9      ====        add a1, s4, s1
                                                  30'd    7625    : data = 32'h    41BF50B3    ;    //    sra x1 x30 x27      ====        sra ra, t5, s11
                                                  30'd    7626    : data = 32'h    CEE1C013    ;    //    xori x0 x3 -786      ====        xori zero, gp, -786
                                                  30'd    7627    : data = 32'h    C0270D13    ;    //    addi x26 x14 -1022      ====        addi s10, a4, -1022
                                                  30'd    7628    : data = 32'h    FA308993    ;    //    addi x19 x1 -93      ====        addi s3, ra, -93
                                                  30'd    7629    : data = 32'h    00575993    ;    //    srli x19 x14 5      ====        srli s3, a4, 5
                                                  30'd    7630    : data = 32'h    01891193    ;    //    slli x3 x18 24      ====        slli gp, s2, 24
                                                  30'd    7631    : data = 32'h    01FC1193    ;    //    slli x3 x24 31      ====        slli gp, s8, 31
                                                  30'd    7632    : data = 32'h    01D38133    ;    //    add x2 x7 x29      ====        add sp, t2, t4
                                                  30'd    7633    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7634    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7635    : data = 32'h    002B30B3    ;    //    sltu x1 x22 x2      ====        sltu ra, s6, sp
                                                  30'd    7636    : data = 32'h    00AFF4B3    ;    //    and x9 x31 x10      ====        and s1, t6, a0
                                                  30'd    7637    : data = 32'h    01231713    ;    //    slli x14 x6 18      ====        slli a4, t1, 18
                                                  30'd    7638    : data = 32'h    40315FB3    ;    //    sra x31 x2 x3      ====        sra t6, sp, gp
                                                  30'd    7639    : data = 32'h    015E0633    ;    //    add x12 x28 x21      ====        add a2, t3, s5
                                                  30'd    7640    : data = 32'h    01E2B0B3    ;    //    sltu x1 x5 x30      ====        sltu ra, t0, t5
                                                  30'd    7641    : data = 32'h    418D8EB3    ;    //    sub x29 x27 x24      ====        sub t4, s11, s8
                                                  30'd    7642    : data = 32'h    01BDBAB3    ;    //    sltu x21 x27 x27      ====        sltu s5, s11, s11
                                                  30'd    7643    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7644    : data = 32'h    ADEC4797    ;    //    auipc x15 712388      ====        auipc a5, 712388
                                                  30'd    7645    : data = 32'h    E423C293    ;    //    xori x5 x7 -446      ====        xori t0, t2, -446
                                                  30'd    7646    : data = 32'h    0085E1B3    ;    //    or x3 x11 x8      ====        or gp, a1, s0
                                                  30'd    7647    : data = 32'h    006F95B3    ;    //    sll x11 x31 x6      ====        sll a1, t6, t1
                                                  30'd    7648    : data = 32'h    01210133    ;    //    add x2 x2 x18      ====        add sp, sp, s2
                                                  30'd    7649    : data = 32'h    40685133    ;    //    sra x2 x16 x6      ====        sra sp, a6, t1
                                                  30'd    7650    : data = 32'h    40608D33    ;    //    sub x26 x1 x6      ====        sub s10, ra, t1
                                                  30'd    7651    : data = 32'h    01810A33    ;    //    add x20 x2 x24      ====        add s4, sp, s8
                                                  30'd    7652    : data = 32'h    D6B7E413    ;    //    ori x8 x15 -661      ====        ori s0, a5, -661
                                                  30'd    7653    : data = 32'h    A27AA013    ;    //    slti x0 x21 -1497      ====        slti zero, s5, -1497
                                                  30'd    7654    : data = 32'h    022873B7    ;    //    lui x7 8839      ====        lui t2, 8839
                                                  30'd    7655    : data = 32'h    342FA093    ;    //    slti x1 x31 834      ====        slti ra, t6, 834
                                                  30'd    7656    : data = 32'h    009921B3    ;    //    slt x3 x18 x9      ====        slt gp, s2, s1
                                                  30'd    7657    : data = 32'h    01E7B6B3    ;    //    sltu x13 x15 x30      ====        sltu a3, a5, t5
                                                  30'd    7658    : data = 32'h    00528C33    ;    //    add x24 x5 x5      ====        add s8, t0, t0
                                                  30'd    7659    : data = 32'h    40B55613    ;    //    srai x12 x10 11      ====        srai a2, a0, 11
                                                  30'd    7660    : data = 32'h    29102617    ;    //    auipc x12 168194      ====        auipc a2, 168194
                                                  30'd    7661    : data = 32'h    00E1D7B3    ;    //    srl x15 x3 x14      ====        srl a5, gp, a4
                                                  30'd    7662    : data = 32'h    0119C4B3    ;    //    xor x9 x19 x17      ====        xor s1, s3, a7
                                                  30'd    7663    : data = 32'h    40E85D33    ;    //    sra x26 x16 x14      ====        sra s10, a6, a4
                                                  30'd    7664    : data = 32'h    012D9D13    ;    //    slli x26 x27 18      ====        slli s10, s11, 18
                                                  30'd    7665    : data = 32'h    01C68633    ;    //    add x12 x13 x28      ====        add a2, a3, t3
                                                  30'd    7666    : data = 32'h    DF058C93    ;    //    addi x25 x11 -528      ====        addi s9, a1, -528
                                                  30'd    7667    : data = 32'h    002C6033    ;    //    or x0 x24 x2      ====        or zero, s8, sp
                                                  30'd    7668    : data = 32'h    DF744617    ;    //    auipc x12 915268      ====        auipc a2, 915268
                                                  30'd    7669    : data = 32'h    00A0F9B3    ;    //    and x19 x1 x10      ====        and s3, ra, a0
                                                  30'd    7670    : data = 32'h    01142133    ;    //    slt x2 x8 x17      ====        slt sp, s0, a7
                                                  30'd    7671    : data = 32'h    40E8D333    ;    //    sra x6 x17 x14      ====        sra t1, a7, a4
                                                  30'd    7672    : data = 32'h    B9DB8413    ;    //    addi x8 x23 -1123      ====        addi s0, s7, -1123
                                                  30'd    7673    : data = 32'h    00BA9433    ;    //    sll x8 x21 x11      ====        sll s0, s5, a1
                                                  30'd    7674    : data = 32'h    00F167B3    ;    //    or x15 x2 x15      ====        or a5, sp, a5
                                                  30'd    7675    : data = 32'h    001B1B33    ;    //    sll x22 x22 x1      ====        sll s6, s6, ra
                                                  30'd    7676    : data = 32'h    41A55D33    ;    //    sra x26 x10 x26      ====        sra s10, a0, s10
                                                  30'd    7677    : data = 32'h    FE5F8193    ;    //    addi x3 x31 -27      ====        addi gp, t6, -27
                                                  30'd    7678    : data = 32'h    F6C74193    ;    //    xori x3 x14 -148      ====        xori gp, a4, -148
                                                  30'd    7679    : data = 32'h    000732B3    ;    //    sltu x5 x14 x0      ====        sltu t0, a4, zero
                                                  30'd    7680    : data = 32'h    4069DC13    ;    //    srai x24 x19 6      ====        srai s8, s3, 6
                                                  30'd    7681    : data = 32'h    0106EA33    ;    //    or x20 x13 x16      ====        or s4, a3, a6
                                                  30'd    7682    : data = 32'h    41085033    ;    //    sra x0 x16 x16      ====        sra zero, a6, a6
                                                  30'd    7683    : data = 32'h    01865333    ;    //    srl x6 x12 x24      ====        srl t1, a2, s8
                                                  30'd    7684    : data = 32'h    005FFFB3    ;    //    and x31 x31 x5      ====        and t6, t6, t0
                                                  30'd    7685    : data = 32'h    00785713    ;    //    srli x14 x16 7      ====        srli a4, a6, 7
                                                  30'd    7686    : data = 32'h    18463097    ;    //    auipc x1 99427      ====        auipc ra, 99427
                                                  30'd    7687    : data = 32'h    414C8C33    ;    //    sub x24 x25 x20      ====        sub s8, s9, s4
                                                  30'd    7688    : data = 32'h    679A7813    ;    //    andi x16 x20 1657      ====        andi a6, s4, 1657
                                                  30'd    7689    : data = 32'h    00A8B5B3    ;    //    sltu x11 x17 x10      ====        sltu a1, a7, a0
                                                  30'd    7690    : data = 32'h    41B8DA33    ;    //    sra x20 x17 x27      ====        sra s4, a7, s11
                                                  30'd    7691    : data = 32'h    53917E93    ;    //    andi x29 x2 1337      ====        andi t4, sp, 1337
                                                  30'd    7692    : data = 32'h    0037ACB3    ;    //    slt x25 x15 x3      ====        slt s9, a5, gp
                                                  30'd    7693    : data = 32'h    00393B33    ;    //    sltu x22 x18 x3      ====        sltu s6, s2, gp
                                                  30'd    7694    : data = 32'h    00ACD6B3    ;    //    srl x13 x25 x10      ====        srl a3, s9, a0
                                                  30'd    7695    : data = 32'h    B0566713    ;    //    ori x14 x12 -1275      ====        ori a4, a2, -1275
                                                  30'd    7696    : data = 32'h    72CC8893    ;    //    addi x17 x25 1836      ====        addi a7, s9, 1836
                                                  30'd    7697    : data = 32'h    01D5DA13    ;    //    srli x20 x11 29      ====        srli s4, a1, 29
                                                  30'd    7698    : data = 32'h    5501C893    ;    //    xori x17 x3 1360      ====        xori a7, gp, 1360
                                                  30'd    7699    : data = 32'h    7080E413    ;    //    ori x8 x1 1800      ====        ori s0, ra, 1800
                                                  30'd    7700    : data = 32'h    3696CD13    ;    //    xori x26 x13 873      ====        xori s10, a3, 873
                                                  30'd    7701    : data = 32'h    0023E1B3    ;    //    or x3 x7 x2      ====        or gp, t2, sp
                                                  30'd    7702    : data = 32'h    EC47F013    ;    //    andi x0 x15 -316      ====        andi zero, a5, -316
                                                  30'd    7703    : data = 32'h    FC22B313    ;    //    sltiu x6 x5 -62      ====        sltiu t1, t0, -62
                                                  30'd    7704    : data = 32'h    01B1AC33    ;    //    slt x24 x3 x27      ====        slt s8, gp, s11
                                                  30'd    7705    : data = 32'h    11286713    ;    //    ori x14 x16 274      ====        ori a4, a6, 274
                                                  30'd    7706    : data = 32'h    003F3733    ;    //    sltu x14 x30 x3      ====        sltu a4, t5, gp
                                                  30'd    7707    : data = 32'h    00071B13    ;    //    slli x22 x14 0      ====        slli s6, a4, 0
                                                  30'd    7708    : data = 32'h    B3773893    ;    //    sltiu x17 x14 -1225      ====        sltiu a7, a4, -1225
                                                  30'd    7709    : data = 32'h    00B85D33    ;    //    srl x26 x16 x11      ====        srl s10, a6, a1
                                                  30'd    7710    : data = 32'h    015364B3    ;    //    or x9 x6 x21      ====        or s1, t1, s5
                                                  30'd    7711    : data = 32'h    4069DF93    ;    //    srai x31 x19 6      ====        srai t6, s3, 6
                                                  30'd    7712    : data = 32'h    628F0F93    ;    //    addi x31 x30 1576      ====        addi t6, t5, 1576
                                                  30'd    7713    : data = 32'h    32477613    ;    //    andi x12 x14 804      ====        andi a2, a4, 804
                                                  30'd    7714    : data = 32'h    E8E36F93    ;    //    ori x31 x6 -370      ====        ori t6, t1, -370
                                                  30'd    7715    : data = 32'h    01782433    ;    //    slt x8 x16 x23      ====        slt s0, a6, s7
                                                  30'd    7716    : data = 32'h    AD034713    ;    //    xori x14 x6 -1328      ====        xori a4, t1, -1328
                                                  30'd    7717    : data = 32'h    9B667993    ;    //    andi x19 x12 -1610      ====        andi s3, a2, -1610
                                                  30'd    7718    : data = 32'h    BE3DE913    ;    //    ori x18 x27 -1053      ====        ori s2, s11, -1053
                                                  30'd    7719    : data = 32'h    0071B033    ;    //    sltu x0 x3 x7      ====        sltu zero, gp, t2
                                                  30'd    7720    : data = 32'h    00216D33    ;    //    or x26 x2 x2      ====        or s10, sp, sp
                                                  30'd    7721    : data = 32'h    59450B13    ;    //    addi x22 x10 1428      ====        addi s6, a0, 1428
                                                  30'd    7722    : data = 32'h    9173E413    ;    //    ori x8 x7 -1769      ====        ori s0, t2, -1769
                                                  30'd    7723    : data = 32'h    000CD8B3    ;    //    srl x17 x25 x0      ====        srl a7, s9, zero
                                                  30'd    7724    : data = 32'h    EA0A7893    ;    //    andi x17 x20 -352      ====        andi a7, s4, -352
                                                  30'd    7725    : data = 32'h    01B98933    ;    //    add x18 x19 x27      ====        add s2, s3, s11
                                                  30'd    7726    : data = 32'h    0104CA33    ;    //    xor x20 x9 x16      ====        xor s4, s1, a6
                                                  30'd    7727    : data = 32'h    1544F193    ;    //    andi x3 x9 340      ====        andi gp, s1, 340
                                                  30'd    7728    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7729    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7730    : data = 32'h    01555833    ;    //    srl x16 x10 x21      ====        srl a6, a0, s5
                                                  30'd    7731    : data = 32'h    B9CEFE17    ;    //    auipc x28 761071      ====        auipc t3, 761071
                                                  30'd    7732    : data = 32'h    0100F2B3    ;    //    and x5 x1 x16      ====        and t0, ra, a6
                                                  30'd    7733    : data = 32'h    0118DAB3    ;    //    srl x21 x17 x17      ====        srl s5, a7, a7
                                                  30'd    7734    : data = 32'h    3B44B813    ;    //    sltiu x16 x9 948      ====        sltiu a6, s1, 948
                                                  30'd    7735    : data = 32'h    A42F0413    ;    //    addi x8 x30 -1470      ====        addi s0, t5, -1470
                                                  30'd    7736    : data = 32'h    49FEF313    ;    //    andi x6 x29 1183      ====        andi t1, t4, 1183
                                                  30'd    7737    : data = 32'h    00D50E33    ;    //    add x28 x10 x13      ====        add t3, a0, a3
                                                  30'd    7738    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7739    : data = 32'h    41F7DF93    ;    //    srai x31 x15 31      ====        srai t6, a5, 31
                                                  30'd    7740    : data = 32'h    6DF7F713    ;    //    andi x14 x15 1759      ====        andi a4, a5, 1759
                                                  30'd    7741    : data = 32'h    41F0DA93    ;    //    srai x21 x1 31      ====        srai s5, ra, 31
                                                  30'd    7742    : data = 32'h    01792933    ;    //    slt x18 x18 x23      ====        slt s2, s2, s7
                                                  30'd    7743    : data = 32'h    00A164B3    ;    //    or x9 x2 x10      ====        or s1, sp, a0
                                                  30'd    7744    : data = 32'h    7D900593    ;    //    addi x11 x0 2009      ====        addi a1, zero, 2009
                                                  30'd    7745    : data = 32'h    8C42EB13    ;    //    ori x22 x5 -1852      ====        ori s6, t0, -1852
                                                  30'd    7746    : data = 32'h    01685D13    ;    //    srli x26 x16 22      ====        srli s10, a6, 22
                                                  30'd    7747    : data = 32'h    E6EC4193    ;    //    xori x3 x24 -402      ====        xori gp, s8, -402
                                                  30'd    7748    : data = 32'h    662AF293    ;    //    andi x5 x21 1634      ====        andi t0, s5, 1634
                                                  30'd    7749    : data = 32'h    40DBD993    ;    //    srai x19 x23 13      ====        srai s3, s7, 13
                                                  30'd    7750    : data = 32'h    00021193    ;    //    slli x3 x4 0      ====        slli gp, tp, 0
                                                  30'd    7751    : data = 32'h    CB4EF9B7    ;    //    lui x19 832751      ====        lui s3, 832751
                                                  30'd    7752    : data = 32'h    AFE27E93    ;    //    andi x29 x4 -1282      ====        andi t4, tp, -1282
                                                  30'd    7753    : data = 32'h    3C7AFA13    ;    //    andi x20 x21 967      ====        andi s4, s5, 967
                                                  30'd    7754    : data = 32'h    00F6A333    ;    //    slt x6 x13 x15      ====        slt t1, a3, a5
                                                  30'd    7755    : data = 32'h    00BA5B13    ;    //    srli x22 x20 11      ====        srli s6, s4, 11
                                                  30'd    7756    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7757    : data = 32'h    0D95FFB7    ;    //    lui x31 55647      ====        lui t6, 55647
                                                  30'd    7758    : data = 32'h    00E3CAB3    ;    //    xor x21 x7 x14      ====        xor s5, t2, a4
                                                  30'd    7759    : data = 32'h    A320ED13    ;    //    ori x26 x1 -1486      ====        ori s10, ra, -1486
                                                  30'd    7760    : data = 32'h    F9A76997    ;    //    auipc x19 1022582      ====        auipc s3, 1022582
                                                  30'd    7761    : data = 32'h    014D8EB3    ;    //    add x29 x27 x20      ====        add t4, s11, s4
                                                  30'd    7762    : data = 32'h    00FEC2B3    ;    //    xor x5 x29 x15      ====        xor t0, t4, a5
                                                  30'd    7763    : data = 32'h    00C285B3    ;    //    add x11 x5 x12      ====        add a1, t0, a2
                                                  30'd    7764    : data = 32'h    7A9C4D93    ;    //    xori x27 x24 1961      ====        xori s11, s8, 1961
                                                  30'd    7765    : data = 32'h    013D86B3    ;    //    add x13 x27 x19      ====        add a3, s11, s3
                                                  30'd    7766    : data = 32'h    E1F27613    ;    //    andi x12 x4 -481      ====        andi a2, tp, -481
                                                  30'd    7767    : data = 32'h    B70E2A13    ;    //    slti x20 x28 -1168      ====        slti s4, t3, -1168
                                                  30'd    7768    : data = 32'h    D2A7B693    ;    //    sltiu x13 x15 -726      ====        sltiu a3, a5, -726
                                                  30'd    7769    : data = 32'h    97A18C93    ;    //    addi x25 x3 -1670      ====        addi s9, gp, -1670
                                                  30'd    7770    : data = 32'h    00ECB7B3    ;    //    sltu x15 x25 x14      ====        sltu a5, s9, a4
                                                  30'd    7771    : data = 32'h    A24AA093    ;    //    slti x1 x21 -1500      ====        slti ra, s5, -1500
                                                  30'd    7772    : data = 32'h    45587013    ;    //    andi x0 x16 1109      ====        andi zero, a6, 1109
                                                  30'd    7773    : data = 32'h    015C4633    ;    //    xor x12 x24 x21      ====        xor a2, s8, s5
                                                  30'd    7774    : data = 32'h    000BA733    ;    //    slt x14 x23 x0      ====        slt a4, s7, zero
                                                  30'd    7775    : data = 32'h    60544B13    ;    //    xori x22 x8 1541      ====        xori s6, s0, 1541
                                                  30'd    7776    : data = 32'h    404CD713    ;    //    srai x14 x25 4      ====        srai a4, s9, 4
                                                  30'd    7777    : data = 32'h    00813033    ;    //    sltu x0 x2 x8      ====        sltu zero, sp, s0
                                                  30'd    7778    : data = 32'h    11FDEE13    ;    //    ori x28 x27 287      ====        ori t3, s11, 287
                                                  30'd    7779    : data = 32'h    4A592413    ;    //    slti x8 x18 1189      ====        slti s0, s2, 1189
                                                  30'd    7780    : data = 32'h    00D8CB33    ;    //    xor x22 x17 x13      ====        xor s6, a7, a3
                                                  30'd    7781    : data = 32'h    01F6DD93    ;    //    srli x27 x13 31      ====        srli s11, a3, 31
                                                  30'd    7782    : data = 32'h    89737117    ;    //    auipc x2 562999      ====        auipc sp, 562999
                                                  30'd    7783    : data = 32'h    16D692B7    ;    //    lui x5 93545      ====        lui t0, 93545
                                                  30'd    7784    : data = 32'h    41A35893    ;    //    srai x17 x6 26      ====        srai a7, t1, 26
                                                  30'd    7785    : data = 32'h    9DD88117    ;    //    auipc x2 646536      ====        auipc sp, 646536
                                                  30'd    7786    : data = 32'h    0050CE33    ;    //    xor x28 x1 x5      ====        xor t3, ra, t0
                                                  30'd    7787    : data = 32'h    401E5893    ;    //    srai x17 x28 1      ====        srai a7, t3, 1
                                                  30'd    7788    : data = 32'h    00281413    ;    //    slli x8 x16 2      ====        slli s0, a6, 2
                                                  30'd    7789    : data = 32'h    007E4893    ;    //    xori x17 x28 7      ====        xori a7, t3, 7
                                                  30'd    7790    : data = 32'h    010A2BB3    ;    //    slt x23 x20 x16      ====        slt s7, s4, a6
                                                  30'd    7791    : data = 32'h    01ADD6B3    ;    //    srl x13 x27 x26      ====        srl a3, s11, s10
                                                  30'd    7792    : data = 32'h    00980633    ;    //    add x12 x16 x9      ====        add a2, a6, s1
                                                  30'd    7793    : data = 32'h    00E509B3    ;    //    add x19 x10 x14      ====        add s3, a0, a4
                                                  30'd    7794    : data = 32'h    405D5913    ;    //    srai x18 x26 5      ====        srai s2, s10, 5
                                                  30'd    7795    : data = 32'h    6CC79797    ;    //    auipc x15 445561      ====        auipc a5, 445561
                                                  30'd    7796    : data = 32'h    91490317    ;    //    auipc x6 595088      ====        auipc t1, 595088
                                                  30'd    7797    : data = 32'h    00DF7133    ;    //    and x2 x30 x13      ====        and sp, t5, a3
                                                  30'd    7798    : data = 32'h    01FFE433    ;    //    or x8 x31 x31      ====        or s0, t6, t6
                                                  30'd    7799    : data = 32'h    41E78CB3    ;    //    sub x25 x15 x30      ====        sub s9, a5, t5
                                                  30'd    7800    : data = 32'h    AABB9097    ;    //    auipc x1 699321      ====        auipc ra, 699321
                                                  30'd    7801    : data = 32'h    43320B13    ;    //    addi x22 x4 1075      ====        addi s6, tp, 1075
                                                  30'd    7802    : data = 32'h    01DA9013    ;    //    slli x0 x21 29      ====        slli zero, s5, 29
                                                  30'd    7803    : data = 32'h    5BBEA093    ;    //    slti x1 x29 1467      ====        slti ra, t4, 1467
                                                  30'd    7804    : data = 32'h    01698733    ;    //    add x14 x19 x22      ====        add a4, s3, s6
                                                  30'd    7805    : data = 32'h    01511FB3    ;    //    sll x31 x2 x21      ====        sll t6, sp, s5
                                                  30'd    7806    : data = 32'h    00006133    ;    //    or x2 x0 x0      ====        or sp, zero, zero
                                                  30'd    7807    : data = 32'h    3844B013    ;    //    sltiu x0 x9 900      ====        sltiu zero, s1, 900
                                                  30'd    7808    : data = 32'h    BACB0593    ;    //    addi x11 x22 -1108      ====        addi a1, s6, -1108
                                                  30'd    7809    : data = 32'h    00F7A733    ;    //    slt x14 x15 x15      ====        slt a4, a5, a5
                                                  30'd    7810    : data = 32'h    392BFB13    ;    //    andi x22 x23 914      ====        andi s6, s7, 914
                                                  30'd    7811    : data = 32'h    E766B837    ;    //    lui x16 947819      ====        lui a6, 947819
                                                  30'd    7812    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7813    : data = 32'h    00A21793    ;    //    slli x15 x4 10      ====        slli a5, tp, 10
                                                  30'd    7814    : data = 32'h    0076FA33    ;    //    and x20 x13 x7      ====        and s4, a3, t2
                                                  30'd    7815    : data = 32'h    00D49F93    ;    //    slli x31 x9 13      ====        slli t6, s1, 13
                                                  30'd    7816    : data = 32'h    00A6D5B3    ;    //    srl x11 x13 x10      ====        srl a1, a3, a0
                                                  30'd    7817    : data = 32'h    AA23C4B7    ;    //    lui x9 696892      ====        lui s1, 696892
                                                  30'd    7818    : data = 32'h    4181D793    ;    //    srai x15 x3 24      ====        srai a5, gp, 24
                                                  30'd    7819    : data = 32'h    00978BB3    ;    //    add x23 x15 x9      ====        add s7, a5, s1
                                                  30'd    7820    : data = 32'h    CDBD2AB7    ;    //    lui x21 842706      ====        lui s5, 842706
                                                  30'd    7821    : data = 32'h    39353D93    ;    //    sltiu x27 x10 915      ====        sltiu s11, a0, 915
                                                  30'd    7822    : data = 32'h    41725C13    ;    //    srai x24 x4 23      ====        srai s8, tp, 23
                                                  30'd    7823    : data = 32'h    88312D93    ;    //    slti x27 x2 -1917      ====        slti s11, sp, -1917
                                                  30'd    7824    : data = 32'h    009ED033    ;    //    srl x0 x29 x9      ====        srl zero, t4, s1
                                                  30'd    7825    : data = 32'h    0B5CE413    ;    //    ori x8 x25 181      ====        ori s0, s9, 181
                                                  30'd    7826    : data = 32'h    01FEC033    ;    //    xor x0 x29 x31      ====        xor zero, t4, t6
                                                  30'd    7827    : data = 32'h    0CA26297    ;    //    auipc x5 51750      ====        auipc t0, 51750
                                                  30'd    7828    : data = 32'h    F57CFE93    ;    //    andi x29 x25 -169      ====        andi t4, s9, -169
                                                  30'd    7829    : data = 32'h    874B4B13    ;    //    xori x22 x22 -1932      ====        xori s6, s6, -1932
                                                  30'd    7830    : data = 32'h    7F93C493    ;    //    xori x9 x7 2041      ====        xori s1, t2, 2041
                                                  30'd    7831    : data = 32'h    000E46B3    ;    //    xor x13 x28 x0      ====        xor a3, t3, zero
                                                  30'd    7832    : data = 32'h    0311AD13    ;    //    slti x26 x3 49      ====        slti s10, gp, 49
                                                  30'd    7833    : data = 32'h    01FD43B3    ;    //    xor x7 x26 x31      ====        xor t2, s10, t6
                                                  30'd    7834    : data = 32'h    007F1633    ;    //    sll x12 x30 x7      ====        sll a2, t5, t2
                                                  30'd    7835    : data = 32'h    00B6D4B3    ;    //    srl x9 x13 x11      ====        srl s1, a3, a1
                                                  30'd    7836    : data = 32'h    40FB5413    ;    //    srai x8 x22 15      ====        srai s0, s6, 15
                                                  30'd    7837    : data = 32'h    004DBFB3    ;    //    sltu x31 x27 x4      ====        sltu t6, s11, tp
                                                  30'd    7838    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7839    : data = 32'h    00E34A33    ;    //    xor x20 x6 x14      ====        xor s4, t1, a4
                                                  30'd    7840    : data = 32'h    008BCDB3    ;    //    xor x27 x23 x8      ====        xor s11, s7, s0
                                                  30'd    7841    : data = 32'h    41B8D5B3    ;    //    sra x11 x17 x27      ====        sra a1, a7, s11
                                                  30'd    7842    : data = 32'h    01313A33    ;    //    sltu x20 x2 x19      ====        sltu s4, sp, s3
                                                  30'd    7843    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7844    : data = 32'h    0044A0B3    ;    //    slt x1 x9 x4      ====        slt ra, s1, tp
                                                  30'd    7845    : data = 32'h    41380433    ;    //    sub x8 x16 x19      ====        sub s0, a6, s3
                                                  30'd    7846    : data = 32'h    41B400B3    ;    //    sub x1 x8 x27      ====        sub ra, s0, s11
                                                  30'd    7847    : data = 32'h    C6097D13    ;    //    andi x26 x18 -928      ====        andi s10, s2, -928
                                                  30'd    7848    : data = 32'h    00345FB3    ;    //    srl x31 x8 x3      ====        srl t6, s0, gp
                                                  30'd    7849    : data = 32'h    00C14833    ;    //    xor x16 x2 x12      ====        xor a6, sp, a2
                                                  30'd    7850    : data = 32'h    406C8833    ;    //    sub x16 x25 x6      ====        sub a6, s9, t1
                                                  30'd    7851    : data = 32'h    7E464A13    ;    //    xori x20 x12 2020      ====        xori s4, a2, 2020
                                                  30'd    7852    : data = 32'h    018036B3    ;    //    sltu x13 x0 x24      ====        sltu a3, zero, s8
                                                  30'd    7853    : data = 32'h    DEB1E817    ;    //    auipc x16 912158      ====        auipc a6, 912158
                                                  30'd    7854    : data = 32'h    3A8533B7    ;    //    lui x7 239699      ====        lui t2, 239699
                                                  30'd    7855    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7856    : data = 32'h    75B13C13    ;    //    sltiu x24 x2 1883      ====        sltiu s8, sp, 1883
                                                  30'd    7857    : data = 32'h    0150D693    ;    //    srli x13 x1 21      ====        srli a3, ra, 21
                                                  30'd    7858    : data = 32'h    AC4EDD17    ;    //    auipc x26 705773      ====        auipc s10, 705773
                                                  30'd    7859    : data = 32'h    631CF013    ;    //    andi x0 x25 1585      ====        andi zero, s9, 1585
                                                  30'd    7860    : data = 32'h    011C5B13    ;    //    srli x22 x24 17      ====        srli s6, s8, 17
                                                  30'd    7861    : data = 32'h    016B29B3    ;    //    slt x19 x22 x22      ====        slt s3, s6, s6
                                                  30'd    7862    : data = 32'h    419B5633    ;    //    sra x12 x22 x25      ====        sra a2, s6, s9
                                                  30'd    7863    : data = 32'h    001EA633    ;    //    slt x12 x29 x1      ====        slt a2, t4, ra
                                                  30'd    7864    : data = 32'h    01C64E33    ;    //    xor x28 x12 x28      ====        xor t3, a2, t3
                                                  30'd    7865    : data = 32'h    01037D33    ;    //    and x26 x6 x16      ====        and s10, t1, a6
                                                  30'd    7866    : data = 32'h    01667FB3    ;    //    and x31 x12 x22      ====        and t6, a2, s6
                                                  30'd    7867    : data = 32'h    69620A93    ;    //    addi x21 x4 1686      ====        addi s5, tp, 1686
                                                  30'd    7868    : data = 32'h    79BFDC37    ;    //    lui x24 498685      ====        lui s8, 498685
                                                  30'd    7869    : data = 32'h    E1868437    ;    //    lui x8 923752      ====        lui s0, 923752
                                                  30'd    7870    : data = 32'h    24DF6193    ;    //    ori x3 x30 589      ====        ori gp, t5, 589
                                                  30'd    7871    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7872    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7873    : data = 32'h    15814713    ;    //    xori x14 x2 344      ====        xori a4, sp, 344
                                                  30'd    7874    : data = 32'h    00BEB393    ;    //    sltiu x7 x29 11      ====        sltiu t2, t4, 11
                                                  30'd    7875    : data = 32'h    01AFE733    ;    //    or x14 x31 x26      ====        or a4, t6, s10
                                                  30'd    7876    : data = 32'h    0178F2B3    ;    //    and x5 x17 x23      ====        and t0, a7, s7
                                                  30'd    7877    : data = 32'h    0176A633    ;    //    slt x12 x13 x23      ====        slt a2, a3, s7
                                                  30'd    7878    : data = 32'h    0160D313    ;    //    srli x6 x1 22      ====        srli t1, ra, 22
                                                  30'd    7879    : data = 32'h    418D8433    ;    //    sub x8 x27 x24      ====        sub s0, s11, s8
                                                  30'd    7880    : data = 32'h    009AE933    ;    //    or x18 x21 x9      ====        or s2, s5, s1
                                                  30'd    7881    : data = 32'h    010CE0B3    ;    //    or x1 x25 x16      ====        or ra, s9, a6
                                                  30'd    7882    : data = 32'h    002B29B3    ;    //    slt x19 x22 x2      ====        slt s3, s6, sp
                                                  30'd    7883    : data = 32'h    C06EA997    ;    //    auipc x19 788202      ====        auipc s3, 788202
                                                  30'd    7884    : data = 32'h    404FDEB3    ;    //    sra x29 x31 x4      ====        sra t4, t6, tp
                                                  30'd    7885    : data = 32'h    015809B3    ;    //    add x19 x16 x21      ====        add s3, a6, s5
                                                  30'd    7886    : data = 32'h    46D76493    ;    //    ori x9 x14 1133      ====        ori s1, a4, 1133
                                                  30'd    7887    : data = 32'h    A21D3B13    ;    //    sltiu x22 x26 -1503      ====        sltiu s6, s10, -1503
                                                  30'd    7888    : data = 32'h    18854A13    ;    //    xori x20 x10 392      ====        xori s4, a0, 392
                                                  30'd    7889    : data = 32'h    AA620713    ;    //    addi x14 x4 -1370      ====        addi a4, tp, -1370
                                                  30'd    7890    : data = 32'h    01BE97B3    ;    //    sll x15 x29 x27      ====        sll a5, t4, s11
                                                  30'd    7891    : data = 32'h    018DDEB3    ;    //    srl x29 x27 x24      ====        srl t4, s11, s8
                                                  30'd    7892    : data = 32'h    6AD5C937    ;    //    lui x18 437596      ====        lui s2, 437596
                                                  30'd    7893    : data = 32'h    005A9E33    ;    //    sll x28 x21 x5      ====        sll t3, s5, t0
                                                  30'd    7894    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7895    : data = 32'h    0107E833    ;    //    or x16 x15 x16      ====        or a6, a5, a6
                                                  30'd    7896    : data = 32'h    01E488B3    ;    //    add x17 x9 x30      ====        add a7, s1, t5
                                                  30'd    7897    : data = 32'h    BB0B0417    ;    //    auipc x8 766128      ====        auipc s0, 766128
                                                  30'd    7898    : data = 32'h    619CDB37    ;    //    lui x22 399821      ====        lui s6, 399821
                                                  30'd    7899    : data = 32'h    00D719B3    ;    //    sll x19 x14 x13      ====        sll s3, a4, a3
                                                  30'd    7900    : data = 32'h    0EFBC0B7    ;    //    lui x1 61372      ====        lui ra, 61372
                                                  30'd    7901    : data = 32'h    CD9A4713    ;    //    xori x14 x20 -807      ====        xori a4, s4, -807
                                                  30'd    7902    : data = 32'h    40A389B3    ;    //    sub x19 x7 x10      ====        sub s3, t2, a0
                                                  30'd    7903    : data = 32'h    40190633    ;    //    sub x12 x18 x1      ====        sub a2, s2, ra
                                                  30'd    7904    : data = 32'h    0061A333    ;    //    slt x6 x3 x6      ====        slt t1, gp, t1
                                                  30'd    7905    : data = 32'h    401D5893    ;    //    srai x17 x26 1      ====        srai a7, s10, 1
                                                  30'd    7906    : data = 32'h    01423B33    ;    //    sltu x22 x4 x20      ====        sltu s6, tp, s4
                                                  30'd    7907    : data = 32'h    00FB5333    ;    //    srl x6 x22 x15      ====        srl t1, s6, a5
                                                  30'd    7908    : data = 32'h    0173BA33    ;    //    sltu x20 x7 x23      ====        sltu s4, t2, s7
                                                  30'd    7909    : data = 32'h    9204B413    ;    //    sltiu x8 x9 -1760      ====        sltiu s0, s1, -1760
                                                  30'd    7910    : data = 32'h    633FAE93    ;    //    slti x29 x31 1587      ====        slti t4, t6, 1587
                                                  30'd    7911    : data = 32'h    89932D13    ;    //    slti x26 x6 -1895      ====        slti s10, t1, -1895
                                                  30'd    7912    : data = 32'h    A1E02793    ;    //    slti x15 x0 -1506      ====        slti a5, zero, -1506
                                                  30'd    7913    : data = 32'h    41FBDC13    ;    //    srai x24 x23 31      ====        srai s8, s7, 31
                                                  30'd    7914    : data = 32'h    FB4D4693    ;    //    xori x13 x26 -76      ====        xori a3, s10, -76
                                                  30'd    7915    : data = 32'h    01E8BFB3    ;    //    sltu x31 x17 x30      ====        sltu t6, a7, t5
                                                  30'd    7916    : data = 32'h    4781A393    ;    //    slti x7 x3 1144      ====        slti t2, gp, 1144
                                                  30'd    7917    : data = 32'h    41025E33    ;    //    sra x28 x4 x16      ====        sra t3, tp, a6
                                                  30'd    7918    : data = 32'h    00FF0433    ;    //    add x8 x30 x15      ====        add s0, t5, a5
                                                  30'd    7919    : data = 32'h    00B25693    ;    //    srli x13 x4 11      ====        srli a3, tp, 11
                                                  30'd    7920    : data = 32'h    00FE3FB3    ;    //    sltu x31 x28 x15      ====        sltu t6, t3, a5
                                                  30'd    7921    : data = 32'h    002BDD13    ;    //    srli x26 x23 2      ====        srli s10, s7, 2
                                                  30'd    7922    : data = 32'h    010A62B3    ;    //    or x5 x20 x16      ====        or t0, s4, a6
                                                  30'd    7923    : data = 32'h    00C32033    ;    //    slt x0 x6 x12      ====        slt zero, t1, a2
                                                  30'd    7924    : data = 32'h    010DAFB3    ;    //    slt x31 x27 x16      ====        slt t6, s11, a6
                                                  30'd    7925    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7926    : data = 32'h    84852793    ;    //    slti x15 x10 -1976      ====        slti a5, a0, -1976
                                                  30'd    7927    : data = 32'h    F7F33D13    ;    //    sltiu x26 x6 -129      ====        sltiu s10, t1, -129
                                                  30'd    7928    : data = 32'h    5D442C93    ;    //    slti x25 x8 1492      ====        slti s9, s0, 1492
                                                  30'd    7929    : data = 32'h    CBAAC037    ;    //    lui x0 834220      ====        lui zero, 834220
                                                  30'd    7930    : data = 32'h    00BD9413    ;    //    slli x8 x27 11      ====        slli s0, s11, 11
                                                  30'd    7931    : data = 32'h    ADE76C93    ;    //    ori x25 x14 -1314      ====        ori s9, a4, -1314
                                                  30'd    7932    : data = 32'h    00BC7133    ;    //    and x2 x24 x11      ====        and sp, s8, a1
                                                  30'd    7933    : data = 32'h    94EE3613    ;    //    sltiu x12 x28 -1714      ====        sltiu a2, t3, -1714
                                                  30'd    7934    : data = 32'h    00C1F633    ;    //    and x12 x3 x12      ====        and a2, gp, a2
                                                  30'd    7935    : data = 32'h    00F18D33    ;    //    add x26 x3 x15      ====        add s10, gp, a5
                                                  30'd    7936    : data = 32'h    00563733    ;    //    sltu x14 x12 x5      ====        sltu a4, a2, t0
                                                  30'd    7937    : data = 32'h    01C29793    ;    //    slli x15 x5 28      ====        slli a5, t0, 28
                                                  30'd    7938    : data = 32'h    FC0A8E13    ;    //    addi x28 x21 -64      ====        addi t3, s5, -64
                                                  30'd    7939    : data = 32'h    001F3833    ;    //    sltu x16 x30 x1      ====        sltu a6, t5, ra
                                                  30'd    7940    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7941    : data = 32'h    016A6633    ;    //    or x12 x20 x22      ====        or a2, s4, s6
                                                  30'd    7942    : data = 32'h    01E3A333    ;    //    slt x6 x7 x30      ====        slt t1, t2, t5
                                                  30'd    7943    : data = 32'h    41B1DFB3    ;    //    sra x31 x3 x27      ====        sra t6, gp, s11
                                                  30'd    7944    : data = 32'h    CA846E93    ;    //    ori x29 x8 -856      ====        ori t4, s0, -856
                                                  30'd    7945    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    7946    : data = 32'h    4F988A13    ;    //    addi x20 x17 1273      ====        addi s4, a7, 1273
                                                  30'd    7947    : data = 32'h    01E19913    ;    //    slli x18 x3 30      ====        slli s2, gp, 30
                                                  30'd    7948    : data = 32'h    01419A13    ;    //    slli x20 x3 20      ====        slli s4, gp, 20
                                                  30'd    7949    : data = 32'h    23979D17    ;    //    auipc x26 145785      ====        auipc s10, 145785
                                                  30'd    7950    : data = 32'h    0093D6B3    ;    //    srl x13 x7 x9      ====        srl a3, t2, s1
                                                  30'd    7951    : data = 32'h    01D4A333    ;    //    slt x6 x9 x29      ====        slt t1, s1, t4
                                                  30'd    7952    : data = 32'h    000E6333    ;    //    or x6 x28 x0      ====        or t1, t3, zero
                                                  30'd    7953    : data = 32'h    4179D633    ;    //    sra x12 x19 x23      ====        sra a2, s3, s7
                                                  30'd    7954    : data = 32'h    40485033    ;    //    sra x0 x16 x4      ====        sra zero, a6, tp
                                                  30'd    7955    : data = 32'h    EE7A4893    ;    //    xori x17 x20 -281      ====        xori a7, s4, -281
                                                  30'd    7956    : data = 32'h    0138FB33    ;    //    and x22 x17 x19      ====        and s6, a7, s3
                                                  30'd    7957    : data = 32'h    001D1333    ;    //    sll x6 x26 x1      ====        sll t1, s10, ra
                                                  30'd    7958    : data = 32'h    0714C837    ;    //    lui x16 29004      ====        lui a6, 29004
                                                  30'd    7959    : data = 32'h    00C75813    ;    //    srli x16 x14 12      ====        srli a6, a4, 12
                                                  30'd    7960    : data = 32'h    4192DD13    ;    //    srai x26 x5 25      ====        srai s10, t0, 25
                                                  30'd    7961    : data = 32'h    0058E3B3    ;    //    or x7 x17 x5      ====        or t2, a7, t0
                                                  30'd    7962    : data = 32'h    41225D93    ;    //    srai x27 x4 18      ====        srai s11, tp, 18
                                                  30'd    7963    : data = 32'h    4EB58E13    ;    //    addi x28 x11 1259      ====        addi t3, a1, 1259
                                                  30'd    7964    : data = 32'h    4007D913    ;    //    srai x18 x15 0      ====        srai s2, a5, 0
                                                  30'd    7965    : data = 32'h    00237B33    ;    //    and x22 x6 x2      ====        and s6, t1, sp
                                                  30'd    7966    : data = 32'h    00B18733    ;    //    add x14 x3 x11      ====        add a4, gp, a1
                                                  30'd    7967    : data = 32'h    01554B33    ;    //    xor x22 x10 x21      ====        xor s6, a0, s5
                                                  30'd    7968    : data = 32'h    57D7F317    ;    //    auipc x6 359807      ====        auipc t1, 359807
                                                  30'd    7969    : data = 32'h    00AF1493    ;    //    slli x9 x30 10      ====        slli s1, t5, 10
                                                  30'd    7970    : data = 32'h    6F534D93    ;    //    xori x27 x6 1781      ====        xori s11, t1, 1781
                                                  30'd    7971    : data = 32'h    01812833    ;    //    slt x16 x2 x24      ====        slt a6, sp, s8
                                                  30'd    7972    : data = 32'h    32C4BD17    ;    //    auipc x26 207947      ====        auipc s10, 207947
                                                  30'd    7973    : data = 32'h    008FD113    ;    //    srli x2 x31 8      ====        srli sp, t6, 8
                                                  30'd    7974    : data = 32'h    018DBEB3    ;    //    sltu x29 x27 x24      ====        sltu t4, s11, s8
                                                  30'd    7975    : data = 32'h    66DAB037    ;    //    lui x0 421291      ====        lui zero, 421291
                                                  30'd    7976    : data = 32'h    00EE49B3    ;    //    xor x19 x28 x14      ====        xor s3, t3, a4
                                                  30'd    7977    : data = 32'h    01859D93    ;    //    slli x27 x11 24      ====        slli s11, a1, 24
                                                  30'd    7978    : data = 32'h    52EC85B7    ;    //    lui x11 339656      ====        lui a1, 339656
                                                  30'd    7979    : data = 32'h    400C00B3    ;    //    sub x1 x24 x0      ====        sub ra, s8, zero
                                                  30'd    7980    : data = 32'h    3AFEF613    ;    //    andi x12 x29 943      ====        andi a2, t4, 943
                                                  30'd    7981    : data = 32'h    DE7CF593    ;    //    andi x11 x25 -537      ====        andi a1, s9, -537
                                                  30'd    7982    : data = 32'h    D717F393    ;    //    andi x7 x15 -655      ====        andi t2, a5, -655
                                                  30'd    7983    : data = 32'h    01B7A8B3    ;    //    slt x17 x15 x27      ====        slt a7, a5, s11
                                                  30'd    7984    : data = 32'h    41634697    ;    //    auipc x13 267828      ====        auipc a3, 267828
                                                  30'd    7985    : data = 32'h    004D72B3    ;    //    and x5 x26 x4      ====        and t0, s10, tp
                                                  30'd    7986    : data = 32'h    41175C13    ;    //    srai x24 x14 17      ====        srai s8, a4, 17
                                                  30'd    7987    : data = 32'h    4CAD6A93    ;    //    ori x21 x26 1226      ====        ori s5, s10, 1226
                                                  30'd    7988    : data = 32'h    837B6193    ;    //    ori x3 x22 -1993      ====        ori gp, s6, -1993
                                                  30'd    7989    : data = 32'h    659E3BB7    ;    //    lui x23 416227      ====        lui s7, 416227
                                                  30'd    7990    : data = 32'h    011EC033    ;    //    xor x0 x29 x17      ====        xor zero, t4, a7
                                                  30'd    7991    : data = 32'h    00B4D8B3    ;    //    srl x17 x9 x11      ====        srl a7, s1, a1
                                                  30'd    7992    : data = 32'h    56C47893    ;    //    andi x17 x8 1388      ====        andi a7, s0, 1388
                                                  30'd    7993    : data = 32'h    004C53B3    ;    //    srl x7 x24 x4      ====        srl t2, s8, tp
                                                  30'd    7994    : data = 32'h    0016EA33    ;    //    or x20 x13 x1      ====        or s4, a3, ra
                                                  30'd    7995    : data = 32'h    00DDD1B3    ;    //    srl x3 x27 x13      ====        srl gp, s11, a3
                                                  30'd    7996    : data = 32'h    40C75E93    ;    //    srai x29 x14 12      ====        srai t4, a4, 12
                                                  30'd    7997    : data = 32'h    40485133    ;    //    sra x2 x16 x4      ====        sra sp, a6, tp
                                                  30'd    7998    : data = 32'h    61950793    ;    //    addi x15 x10 1561      ====        addi a5, a0, 1561
                                                  30'd    7999    : data = 32'h    48438437    ;    //    lui x8 295992      ====        lui s0, 295992
                                                  30'd    8000    : data = 32'h    7A8D7A13    ;    //    andi x20 x26 1960      ====        andi s4, s10, 1960
                                                  30'd    8001    : data = 32'h    31A07813    ;    //    andi x16 x0 794      ====        andi a6, zero, 794
                                                  30'd    8002    : data = 32'h    40860633    ;    //    sub x12 x12 x8      ====        sub a2, a2, s0
                                                  30'd    8003    : data = 32'h    328E2D13    ;    //    slti x26 x28 808      ====        slti s10, t3, 808
                                                  30'd    8004    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8005    : data = 32'h    00F4DCB3    ;    //    srl x25 x9 x15      ====        srl s9, s1, a5
                                                  30'd    8006    : data = 32'h    2CB3E717    ;    //    auipc x14 183102      ====        auipc a4, 183102
                                                  30'd    8007    : data = 32'h    359F7593    ;    //    andi x11 x30 857      ====        andi a1, t5, 857
                                                  30'd    8008    : data = 32'h    0041F4B3    ;    //    and x9 x3 x4      ====        and s1, gp, tp
                                                  30'd    8009    : data = 32'h    F3793D13    ;    //    sltiu x26 x18 -201      ====        sltiu s10, s2, -201
                                                  30'd    8010    : data = 32'h    006F90B3    ;    //    sll x1 x31 x6      ====        sll ra, t6, t1
                                                  30'd    8011    : data = 32'h    30DCFB13    ;    //    andi x22 x25 781      ====        andi s6, s9, 781
                                                  30'd    8012    : data = 32'h    4028D893    ;    //    srai x17 x17 2      ====        srai a7, a7, 2
                                                  30'd    8013    : data = 32'h    00DEC2B3    ;    //    xor x5 x29 x13      ====        xor t0, t4, a3
                                                  30'd    8014    : data = 32'h    75E46093    ;    //    ori x1 x8 1886      ====        ori ra, s0, 1886
                                                  30'd    8015    : data = 32'h    413A5413    ;    //    srai x8 x20 19      ====        srai s0, s4, 19
                                                  30'd    8016    : data = 32'h    015CA8B3    ;    //    slt x17 x25 x21      ====        slt a7, s9, s5
                                                  30'd    8017    : data = 32'h    01598133    ;    //    add x2 x19 x21      ====        add sp, s3, s5
                                                  30'd    8018    : data = 32'h    40455D93    ;    //    srai x27 x10 4      ====        srai s11, a0, 4
                                                  30'd    8019    : data = 32'h    AC65ED93    ;    //    ori x27 x11 -1338      ====        ori s11, a1, -1338
                                                  30'd    8020    : data = 32'h    00D358B3    ;    //    srl x17 x6 x13      ====        srl a7, t1, a3
                                                  30'd    8021    : data = 32'h    4129DB93    ;    //    srai x23 x19 18      ====        srai s7, s3, 18
                                                  30'd    8022    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8023    : data = 32'h    C6B1BF97    ;    //    auipc x31 813851      ====        auipc t6, 813851
                                                  30'd    8024    : data = 32'h    41D6D493    ;    //    srai x9 x13 29      ====        srai s1, a3, 29
                                                  30'd    8025    : data = 32'h    008F5E33    ;    //    srl x28 x30 x8      ====        srl t3, t5, s0
                                                  30'd    8026    : data = 32'h    00C4BAB3    ;    //    sltu x21 x9 x12      ====        sltu s5, s1, a2
                                                  30'd    8027    : data = 32'h    00370933    ;    //    add x18 x14 x3      ====        add s2, a4, gp
                                                  30'd    8028    : data = 32'h    01B3DFB3    ;    //    srl x31 x7 x27      ====        srl t6, t2, s11
                                                  30'd    8029    : data = 32'h    004F6833    ;    //    or x16 x30 x4      ====        or a6, t5, tp
                                                  30'd    8030    : data = 32'h    DEC12B13    ;    //    slti x22 x2 -532      ====        slti s6, sp, -532
                                                  30'd    8031    : data = 32'h    00FF74B3    ;    //    and x9 x30 x15      ====        and s1, t5, a5
                                                  30'd    8032    : data = 32'h    412B5A33    ;    //    sra x20 x22 x18      ====        sra s4, s6, s2
                                                  30'd    8033    : data = 32'h    00B45DB3    ;    //    srl x27 x8 x11      ====        srl s11, s0, a1
                                                  30'd    8034    : data = 32'h    01168BB3    ;    //    add x23 x13 x17      ====        add s7, a3, a7
                                                  30'd    8035    : data = 32'h    536D5717    ;    //    auipc x14 341717      ====        auipc a4, 341717
                                                  30'd    8036    : data = 32'h    0065D6B3    ;    //    srl x13 x11 x6      ====        srl a3, a1, t1
                                                  30'd    8037    : data = 32'h    FE164713    ;    //    xori x14 x12 -31      ====        xori a4, a2, -31
                                                  30'd    8038    : data = 32'h    01FDDE13    ;    //    srli x28 x27 31      ====        srli t3, s11, 31
                                                  30'd    8039    : data = 32'h    007192B3    ;    //    sll x5 x3 x7      ====        sll t0, gp, t2
                                                  30'd    8040    : data = 32'h    000D9633    ;    //    sll x12 x27 x0      ====        sll a2, s11, zero
                                                  30'd    8041    : data = 32'h    57714193    ;    //    xori x3 x2 1399      ====        xori gp, sp, 1399
                                                  30'd    8042    : data = 32'h    0107CA33    ;    //    xor x20 x15 x16      ====        xor s4, a5, a6
                                                  30'd    8043    : data = 32'h    41B95A93    ;    //    srai x21 x18 27      ====        srai s5, s2, 27
                                                  30'd    8044    : data = 32'h    EA095C37    ;    //    lui x24 958613      ====        lui s8, 958613
                                                  30'd    8045    : data = 32'h    405F0FB3    ;    //    sub x31 x30 x5      ====        sub t6, t5, t0
                                                  30'd    8046    : data = 32'h    40185293    ;    //    srai x5 x16 1      ====        srai t0, a6, 1
                                                  30'd    8047    : data = 32'h    403DD813    ;    //    srai x16 x27 3      ====        srai a6, s11, 3
                                                  30'd    8048    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8049    : data = 32'h    00F50B33    ;    //    add x22 x10 x15      ====        add s6, a0, a5
                                                  30'd    8050    : data = 32'h    0087CE33    ;    //    xor x28 x15 x8      ====        xor t3, a5, s0
                                                  30'd    8051    : data = 32'h    97832A93    ;    //    slti x21 x6 -1672      ====        slti s5, t1, -1672
                                                  30'd    8052    : data = 32'h    004880B3    ;    //    add x1 x17 x4      ====        add ra, a7, tp
                                                  30'd    8053    : data = 32'h    0038F2B3    ;    //    and x5 x17 x3      ====        and t0, a7, gp
                                                  30'd    8054    : data = 32'h    4EA5A593    ;    //    slti x11 x11 1258      ====        slti a1, a1, 1258
                                                  30'd    8055    : data = 32'h    54D64313    ;    //    xori x6 x12 1357      ====        xori t1, a2, 1357
                                                  30'd    8056    : data = 32'h    66F1E413    ;    //    ori x8 x3 1647      ====        ori s0, gp, 1647
                                                  30'd    8057    : data = 32'h    030D6293    ;    //    ori x5 x26 48      ====        ori t0, s10, 48
                                                  30'd    8058    : data = 32'h    01E66BB3    ;    //    or x23 x12 x30      ====        or s7, a2, t5
                                                  30'd    8059    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8060    : data = 32'h    68A88437    ;    //    lui x8 428680      ====        lui s0, 428680
                                                  30'd    8061    : data = 32'h    40A75733    ;    //    sra x14 x14 x10      ====        sra a4, a4, a0
                                                  30'd    8062    : data = 32'h    00441733    ;    //    sll x14 x8 x4      ====        sll a4, s0, tp
                                                  30'd    8063    : data = 32'h    018A06B3    ;    //    add x13 x20 x24      ====        add a3, s4, s8
                                                  30'd    8064    : data = 32'h    BF750BB7    ;    //    lui x23 784208      ====        lui s7, 784208
                                                  30'd    8065    : data = 32'h    617FC713    ;    //    xori x14 x31 1559      ====        xori a4, t6, 1559
                                                  30'd    8066    : data = 32'h    4124D033    ;    //    sra x0 x9 x18      ====        sra zero, s1, s2
                                                  30'd    8067    : data = 32'h    703F3D13    ;    //    sltiu x26 x30 1795      ====        sltiu s10, t5, 1795
                                                  30'd    8068    : data = 32'h    414000B3    ;    //    sub x1 x0 x20      ====        sub ra, zero, s4
                                                  30'd    8069    : data = 32'h    A9AD7913    ;    //    andi x18 x26 -1382      ====        andi s2, s10, -1382
                                                  30'd    8070    : data = 32'h    00022E33    ;    //    slt x28 x4 x0      ====        slt t3, tp, zero
                                                  30'd    8071    : data = 32'h    004BE633    ;    //    or x12 x23 x4      ====        or a2, s7, tp
                                                  30'd    8072    : data = 32'h    414A5D13    ;    //    srai x26 x20 20      ====        srai s10, s4, 20
                                                  30'd    8073    : data = 32'h    3A5E3113    ;    //    sltiu x2 x28 933      ====        sltiu sp, t3, 933
                                                  30'd    8074    : data = 32'h    B44EFE93    ;    //    andi x29 x29 -1212      ====        andi t4, t4, -1212
                                                  30'd    8075    : data = 32'h    01702933    ;    //    slt x18 x0 x23      ====        slt s2, zero, s7
                                                  30'd    8076    : data = 32'h    A682FF93    ;    //    andi x31 x5 -1432      ====        andi t6, t0, -1432
                                                  30'd    8077    : data = 32'h    405A0CB3    ;    //    sub x25 x20 x5      ====        sub s9, s4, t0
                                                  30'd    8078    : data = 32'h    962D8E17    ;    //    auipc x28 615128      ====        auipc t3, 615128
                                                  30'd    8079    : data = 32'h    0140D1B3    ;    //    srl x3 x1 x20      ====        srl gp, ra, s4
                                                  30'd    8080    : data = 32'h    01E733B3    ;    //    sltu x7 x14 x30      ====        sltu t2, a4, t5
                                                  30'd    8081    : data = 32'h    01C0A8B3    ;    //    slt x17 x1 x28      ====        slt a7, ra, t3
                                                  30'd    8082    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8083    : data = 32'h    00748733    ;    //    add x14 x9 x7      ====        add a4, s1, t2
                                                  30'd    8084    : data = 32'h    41D25CB3    ;    //    sra x25 x4 x29      ====        sra s9, tp, t4
                                                  30'd    8085    : data = 32'h    017E8433    ;    //    add x8 x29 x23      ====        add s0, t4, s7
                                                  30'd    8086    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8087    : data = 32'h    40DBD613    ;    //    srai x12 x23 13      ====        srai a2, s7, 13
                                                  30'd    8088    : data = 32'h    01D20CB3    ;    //    add x25 x4 x29      ====        add s9, tp, t4
                                                  30'd    8089    : data = 32'h    60FB6A13    ;    //    ori x20 x22 1551      ====        ori s4, s6, 1551
                                                  30'd    8090    : data = 32'h    00769313    ;    //    slli x6 x13 7      ====        slli t1, a3, 7
                                                  30'd    8091    : data = 32'h    418501B3    ;    //    sub x3 x10 x24      ====        sub gp, a0, s8
                                                  30'd    8092    : data = 32'h    AB6EB113    ;    //    sltiu x2 x29 -1354      ====        sltiu sp, t4, -1354
                                                  30'd    8093    : data = 32'h    410459B3    ;    //    sra x19 x8 x16      ====        sra s3, s0, a6
                                                  30'd    8094    : data = 32'h    2A553593    ;    //    sltiu x11 x10 677      ====        sltiu a1, a0, 677
                                                  30'd    8095    : data = 32'h    007E9893    ;    //    slli x17 x29 7      ====        slli a7, t4, 7
                                                  30'd    8096    : data = 32'h    0184C933    ;    //    xor x18 x9 x24      ====        xor s2, s1, s8
                                                  30'd    8097    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8098    : data = 32'h    4130DA93    ;    //    srai x21 x1 19      ====        srai s5, ra, 19
                                                  30'd    8099    : data = 32'h    8BE9B913    ;    //    sltiu x18 x19 -1858      ====        sltiu s2, s3, -1858
                                                  30'd    8100    : data = 32'h    D18F4793    ;    //    xori x15 x30 -744      ====        xori a5, t5, -744
                                                  30'd    8101    : data = 32'h    015AE633    ;    //    or x12 x21 x21      ====        or a2, s5, s5
                                                  30'd    8102    : data = 32'h    0014D2B3    ;    //    srl x5 x9 x1      ====        srl t0, s1, ra
                                                  30'd    8103    : data = 32'h    000385B3    ;    //    add x11 x7 x0      ====        add a1, t2, zero
                                                  30'd    8104    : data = 32'h    4C21DD17    ;    //    auipc x26 311837      ====        auipc s10, 311837
                                                  30'd    8105    : data = 32'h    00A040B3    ;    //    xor x1 x0 x10      ====        xor ra, zero, a0
                                                  30'd    8106    : data = 32'h    3BB7E313    ;    //    ori x6 x15 955      ====        ori t1, a5, 955
                                                  30'd    8107    : data = 32'h    404B04B3    ;    //    sub x9 x22 x4      ====        sub s1, s6, tp
                                                  30'd    8108    : data = 32'h    410A56B3    ;    //    sra x13 x20 x16      ====        sra a3, s4, a6
                                                  30'd    8109    : data = 32'h    0B1ECA93    ;    //    xori x21 x29 177      ====        xori s5, t4, 177
                                                  30'd    8110    : data = 32'h    015F48B3    ;    //    xor x17 x30 x21      ====        xor a7, t5, s5
                                                  30'd    8111    : data = 32'h    40AB5933    ;    //    sra x18 x22 x10      ====        sra s2, s6, a0
                                                  30'd    8112    : data = 32'h    010DFCB3    ;    //    and x25 x27 x16      ====        and s9, s11, a6
                                                  30'd    8113    : data = 32'h    019BF6B3    ;    //    and x13 x23 x25      ====        and a3, s7, s9
                                                  30'd    8114    : data = 32'h    00357133    ;    //    and x2 x10 x3      ====        and sp, a0, gp
                                                  30'd    8115    : data = 32'h    411C0EB3    ;    //    sub x29 x24 x17      ====        sub t4, s8, a7
                                                  30'd    8116    : data = 32'h    690D6713    ;    //    ori x14 x26 1680      ====        ori a4, s10, 1680
                                                  30'd    8117    : data = 32'h    001B5633    ;    //    srl x12 x22 x1      ====        srl a2, s6, ra
                                                  30'd    8118    : data = 32'h    0079B133    ;    //    sltu x2 x19 x7      ====        sltu sp, s3, t2
                                                  30'd    8119    : data = 32'h    6B530B37    ;    //    lui x22 439600      ====        lui s6, 439600
                                                  30'd    8120    : data = 32'h    41ABDB13    ;    //    srai x22 x23 26      ====        srai s6, s7, 26
                                                  30'd    8121    : data = 32'h    01A781B3    ;    //    add x3 x15 x26      ====        add gp, a5, s10
                                                  30'd    8122    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8123    : data = 32'h    AE787F93    ;    //    andi x31 x16 -1305      ====        andi t6, a6, -1305
                                                  30'd    8124    : data = 32'h    00D1DB13    ;    //    srli x22 x3 13      ====        srli s6, gp, 13
                                                  30'd    8125    : data = 32'h    25547A93    ;    //    andi x21 x8 597      ====        andi s5, s0, 597
                                                  30'd    8126    : data = 32'h    00124B33    ;    //    xor x22 x4 x1      ====        xor s6, tp, ra
                                                  30'd    8127    : data = 32'h    0108B133    ;    //    sltu x2 x17 x16      ====        sltu sp, a7, a6
                                                  30'd    8128    : data = 32'h    408E5CB3    ;    //    sra x25 x28 x8      ====        sra s9, t3, s0
                                                  30'd    8129    : data = 32'h    41360B33    ;    //    sub x22 x12 x19      ====        sub s6, a2, s3
                                                  30'd    8130    : data = 32'h    415BE293    ;    //    ori x5 x23 1045      ====        ori t0, s7, 1045
                                                  30'd    8131    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8132    : data = 32'h    656CFB93    ;    //    andi x23 x25 1622      ====        andi s7, s9, 1622
                                                  30'd    8133    : data = 32'h    E50FB3B7    ;    //    lui x7 938235      ====        lui t2, 938235
                                                  30'd    8134    : data = 32'h    00A4D093    ;    //    srli x1 x9 10      ====        srli ra, s1, 10
                                                  30'd    8135    : data = 32'h    7C3F0B13    ;    //    addi x22 x30 1987      ====        addi s6, t5, 1987
                                                  30'd    8136    : data = 32'h    012CBAB3    ;    //    sltu x21 x25 x18      ====        sltu s5, s9, s2
                                                  30'd    8137    : data = 32'h    0AA3EB37    ;    //    lui x22 43582      ====        lui s6, 43582
                                                  30'd    8138    : data = 32'h    41E95413    ;    //    srai x8 x18 30      ====        srai s0, s2, 30
                                                  30'd    8139    : data = 32'h    414401B3    ;    //    sub x3 x8 x20      ====        sub gp, s0, s4
                                                  30'd    8140    : data = 32'h    592CE493    ;    //    ori x9 x25 1426      ====        ori s1, s9, 1426
                                                  30'd    8141    : data = 32'h    40D1DFB3    ;    //    sra x31 x3 x13      ====        sra t6, gp, a3
                                                  30'd    8142    : data = 32'h    14C47293    ;    //    andi x5 x8 332      ====        andi t0, s0, 332
                                                  30'd    8143    : data = 32'h    0098C5B3    ;    //    xor x11 x17 x9      ====        xor a1, a7, s1
                                                  30'd    8144    : data = 32'h    04DA8793    ;    //    addi x15 x21 77      ====        addi a5, s5, 77
                                                  30'd    8145    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8146    : data = 32'h    00A19A13    ;    //    slli x20 x3 10      ====        slli s4, gp, 10
                                                  30'd    8147    : data = 32'h    0025F433    ;    //    and x8 x11 x2      ====        and s0, a1, sp
                                                  30'd    8148    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8149    : data = 32'h    01835CB3    ;    //    srl x25 x6 x24      ====        srl s9, t1, s8
                                                  30'd    8150    : data = 32'h    72A3C697    ;    //    auipc x13 469564      ====        auipc a3, 469564
                                                  30'd    8151    : data = 32'h    501E7493    ;    //    andi x9 x28 1281      ====        andi s1, t3, 1281
                                                  30'd    8152    : data = 32'h    C7E4F593    ;    //    andi x11 x9 -898      ====        andi a1, s1, -898
                                                  30'd    8153    : data = 32'h    00D0CD33    ;    //    xor x26 x1 x13      ====        xor s10, ra, a3
                                                  30'd    8154    : data = 32'h    00645813    ;    //    srli x16 x8 6      ====        srli a6, s0, 6
                                                  30'd    8155    : data = 32'h    FB64E993    ;    //    ori x19 x9 -74      ====        ori s3, s1, -74
                                                  30'd    8156    : data = 32'h    9D338A93    ;    //    addi x21 x7 -1581      ====        addi s5, t2, -1581
                                                  30'd    8157    : data = 32'h    004CABB3    ;    //    slt x23 x25 x4      ====        slt s7, s9, tp
                                                  30'd    8158    : data = 32'h    411A07B3    ;    //    sub x15 x20 x17      ====        sub a5, s4, a7
                                                  30'd    8159    : data = 32'h    48D9A917    ;    //    auipc x18 298394      ====        auipc s2, 298394
                                                  30'd    8160    : data = 32'h    41EF8B33    ;    //    sub x22 x31 x30      ====        sub s6, t6, t5
                                                  30'd    8161    : data = 32'h    00B6C733    ;    //    xor x14 x13 x11      ====        xor a4, a3, a1
                                                  30'd    8162    : data = 32'h    00F5FE33    ;    //    and x28 x11 x15      ====        and t3, a1, a5
                                                  30'd    8163    : data = 32'h    CC702F93    ;    //    slti x31 x0 -825      ====        slti t6, zero, -825
                                                  30'd    8164    : data = 32'h    40205713    ;    //    srai x14 x0 2      ====        srai a4, zero, 2
                                                  30'd    8165    : data = 32'h    72C5F493    ;    //    andi x9 x11 1836      ====        andi s1, a1, 1836
                                                  30'd    8166    : data = 32'h    01BE9633    ;    //    sll x12 x29 x27      ====        sll a2, t4, s11
                                                  30'd    8167    : data = 32'h    0044FFB3    ;    //    and x31 x9 x4      ====        and t6, s1, tp
                                                  30'd    8168    : data = 32'h    0176D633    ;    //    srl x12 x13 x23      ====        srl a2, a3, s7
                                                  30'd    8169    : data = 32'h    0142D913    ;    //    srli x18 x5 20      ====        srli s2, t0, 20
                                                  30'd    8170    : data = 32'h    613C6B13    ;    //    ori x22 x24 1555      ====        ori s6, s8, 1555
                                                  30'd    8171    : data = 32'h    0057D793    ;    //    srli x15 x15 5      ====        srli a5, a5, 5
                                                  30'd    8172    : data = 32'h    00ACAA93    ;    //    slti x21 x25 10      ====        slti s5, s9, 10
                                                  30'd    8173    : data = 32'h    227D0D93    ;    //    addi x27 x26 551      ====        addi s11, s10, 551
                                                  30'd    8174    : data = 32'h    0146BA33    ;    //    sltu x20 x13 x20      ====        sltu s4, a3, s4
                                                  30'd    8175    : data = 32'h    01C66BB3    ;    //    or x23 x12 x28      ====        or s7, a2, t3
                                                  30'd    8176    : data = 32'h    00D81793    ;    //    slli x15 x16 13      ====        slli a5, a6, 13
                                                  30'd    8177    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8178    : data = 32'h    4043D6B3    ;    //    sra x13 x7 x4      ====        sra a3, t2, tp
                                                  30'd    8179    : data = 32'h    004959B3    ;    //    srl x19 x18 x4      ====        srl s3, s2, tp
                                                  30'd    8180    : data = 32'h    019D5893    ;    //    srli x17 x26 25      ====        srli a7, s10, 25
                                                  30'd    8181    : data = 32'h    07A44A13    ;    //    xori x20 x8 122      ====        xori s4, s0, 122
                                                  30'd    8182    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8183    : data = 32'h    935E6C13    ;    //    ori x24 x28 -1739      ====        ori s8, t3, -1739
                                                  30'd    8184    : data = 32'h    40A6D8B3    ;    //    sra x17 x13 x10      ====        sra a7, a3, a0
                                                  30'd    8185    : data = 32'h    01845933    ;    //    srl x18 x8 x24      ====        srl s2, s0, s8
                                                  30'd    8186    : data = 32'h    4761F897    ;    //    auipc x17 292383      ====        auipc a7, 292383
                                                  30'd    8187    : data = 32'h    41CD8733    ;    //    sub x14 x27 x28      ====        sub a4, s11, t3
                                                  30'd    8188    : data = 32'h    01C93FB3    ;    //    sltu x31 x18 x28      ====        sltu t6, s2, t3
                                                  30'd    8189    : data = 32'h    00232733    ;    //    slt x14 x6 x2      ====        slt a4, t1, sp
                                                  30'd    8190    : data = 32'h    032FA737    ;    //    lui x14 13050      ====        lui a4, 13050
                                                  30'd    8191    : data = 32'h    007B71B3    ;    //    and x3 x22 x7      ====        and gp, s6, t2
                                                  30'd    8192    : data = 32'h    0086CC33    ;    //    xor x24 x13 x8      ====        xor s8, a3, s0
                                                  30'd    8193    : data = 32'h    01175D93    ;    //    srli x27 x14 17      ====        srli s11, a4, 17
                                                  30'd    8194    : data = 32'h    4002DA93    ;    //    srai x21 x5 0      ====        srai s5, t0, 0
                                                  30'd    8195    : data = 32'h    01A77C33    ;    //    and x24 x14 x26      ====        and s8, a4, s10
                                                  30'd    8196    : data = 32'h    00CCD3B3    ;    //    srl x7 x25 x12      ====        srl t2, s9, a2
                                                  30'd    8197    : data = 32'h    41045C93    ;    //    srai x25 x8 16      ====        srai s9, s0, 16
                                                  30'd    8198    : data = 32'h    01533133    ;    //    sltu x2 x6 x21      ====        sltu sp, t1, s5
                                                  30'd    8199    : data = 32'h    40095A13    ;    //    srai x20 x18 0      ====        srai s4, s2, 0
                                                  30'd    8200    : data = 32'h    00EDC733    ;    //    xor x14 x27 x14      ====        xor a4, s11, a4
                                                  30'd    8201    : data = 32'h    F44D7413    ;    //    andi x8 x26 -188      ====        andi s0, s10, -188
                                                  30'd    8202    : data = 32'h    404802B3    ;    //    sub x5 x16 x4      ====        sub t0, a6, tp
                                                  30'd    8203    : data = 32'h    C6D8E093    ;    //    ori x1 x17 -915      ====        ori ra, a7, -915
                                                  30'd    8204    : data = 32'h    D6E87A13    ;    //    andi x20 x16 -658      ====        andi s4, a6, -658
                                                  30'd    8205    : data = 32'h    01138833    ;    //    add x16 x7 x17      ====        add a6, t2, a7
                                                  30'd    8206    : data = 32'h    209C4313    ;    //    xori x6 x24 521      ====        xori t1, s8, 521
                                                  30'd    8207    : data = 32'h    009E37B3    ;    //    sltu x15 x28 x9      ====        sltu a5, t3, s1
                                                  30'd    8208    : data = 32'h    11D87D13    ;    //    andi x26 x16 285      ====        andi s10, a6, 285
                                                  30'd    8209    : data = 32'h    011FEEB3    ;    //    or x29 x31 x17      ====        or t4, t6, a7
                                                  30'd    8210    : data = 32'h    C1F73113    ;    //    sltiu x2 x14 -993      ====        sltiu sp, a4, -993
                                                  30'd    8211    : data = 32'h    4080D633    ;    //    sra x12 x1 x8      ====        sra a2, ra, s0
                                                  30'd    8212    : data = 32'h    10D2DA37    ;    //    lui x20 68909      ====        lui s4, 68909
                                                  30'd    8213    : data = 32'h    3C2A2D17    ;    //    auipc x26 246434      ====        auipc s10, 246434
                                                  30'd    8214    : data = 32'h    28BF3B13    ;    //    sltiu x22 x30 651      ====        sltiu s6, t5, 651
                                                  30'd    8215    : data = 32'h    002124B3    ;    //    slt x9 x2 x2      ====        slt s1, sp, sp
                                                  30'd    8216    : data = 32'h    81C20713    ;    //    addi x14 x4 -2020      ====        addi a4, tp, -2020
                                                  30'd    8217    : data = 32'h    018E9413    ;    //    slli x8 x29 24      ====        slli s0, t4, 24
                                                  30'd    8218    : data = 32'h    79E82393    ;    //    slti x7 x16 1950      ====        slti t2, a6, 1950
                                                  30'd    8219    : data = 32'h    7C0BCA13    ;    //    xori x20 x23 1984      ====        xori s4, s7, 1984
                                                  30'd    8220    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8221    : data = 32'h    018A5913    ;    //    srli x18 x20 24      ====        srli s2, s4, 24
                                                  30'd    8222    : data = 32'h    A1B3ABB7    ;    //    lui x23 662330      ====        lui s7, 662330
                                                  30'd    8223    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8224    : data = 32'h    41545A13    ;    //    srai x20 x8 21      ====        srai s4, s0, 21
                                                  30'd    8225    : data = 32'h    01BD56B3    ;    //    srl x13 x26 x27      ====        srl a3, s10, s11
                                                  30'd    8226    : data = 32'h    40DC0D33    ;    //    sub x26 x24 x13      ====        sub s10, s8, a3
                                                  30'd    8227    : data = 32'h    01431133    ;    //    sll x2 x6 x20      ====        sll sp, t1, s4
                                                  30'd    8228    : data = 32'h    453D2697    ;    //    auipc x13 283602      ====        auipc a3, 283602
                                                  30'd    8229    : data = 32'h    01B89C93    ;    //    slli x25 x17 27      ====        slli s9, a7, 27
                                                  30'd    8230    : data = 32'h    417F0933    ;    //    sub x18 x30 x23      ====        sub s2, t5, s7
                                                  30'd    8231    : data = 32'h    01076433    ;    //    or x8 x14 x16      ====        or s0, a4, a6
                                                  30'd    8232    : data = 32'h    065B0793    ;    //    addi x15 x22 101      ====        addi a5, s6, 101
                                                  30'd    8233    : data = 32'h    011A9193    ;    //    slli x3 x21 17      ====        slli gp, s5, 17
                                                  30'd    8234    : data = 32'h    00029293    ;    //    slli x5 x5 0      ====        slli t0, t0, 0
                                                  30'd    8235    : data = 32'h    00F93FB3    ;    //    sltu x31 x18 x15      ====        sltu t6, s2, a5
                                                  30'd    8236    : data = 32'h    018858B3    ;    //    srl x17 x16 x24      ====        srl a7, a6, s8
                                                  30'd    8237    : data = 32'h    40F2D033    ;    //    sra x0 x5 x15      ====        sra zero, t0, a5
                                                  30'd    8238    : data = 32'h    91DE8693    ;    //    addi x13 x29 -1763      ====        addi a3, t4, -1763
                                                  30'd    8239    : data = 32'h    0049E933    ;    //    or x18 x19 x4      ====        or s2, s3, tp
                                                  30'd    8240    : data = 32'h    00E9D393    ;    //    srli x7 x19 14      ====        srli t2, s3, 14
                                                  30'd    8241    : data = 32'h    01991B93    ;    //    slli x23 x18 25      ====        slli s7, s2, 25
                                                  30'd    8242    : data = 32'h    01516333    ;    //    or x6 x2 x21      ====        or t1, sp, s5
                                                  30'd    8243    : data = 32'h    00CE8AB3    ;    //    add x21 x29 x12      ====        add s5, t4, a2
                                                  30'd    8244    : data = 32'h    14B70313    ;    //    addi x6 x14 331      ====        addi t1, a4, 331
                                                  30'd    8245    : data = 32'h    0FECC893    ;    //    xori x17 x25 254      ====        xori a7, s9, 254
                                                  30'd    8246    : data = 32'h    012449B3    ;    //    xor x19 x8 x18      ====        xor s3, s0, s2
                                                  30'd    8247    : data = 32'h    794E0F93    ;    //    addi x31 x28 1940      ====        addi t6, t3, 1940
                                                  30'd    8248    : data = 32'h    0150F2B3    ;    //    and x5 x1 x21      ====        and t0, ra, s5
                                                  30'd    8249    : data = 32'h    86778C17    ;    //    auipc x24 550776      ====        auipc s8, 550776
                                                  30'd    8250    : data = 32'h    01B61033    ;    //    sll x0 x12 x27      ====        sll zero, a2, s11
                                                  30'd    8251    : data = 32'h    1B7FE793    ;    //    ori x15 x31 439      ====        ori a5, t6, 439
                                                  30'd    8252    : data = 32'h    00BF5A33    ;    //    srl x20 x30 x11      ====        srl s4, t5, a1
                                                  30'd    8253    : data = 32'h    4032D933    ;    //    sra x18 x5 x3      ====        sra s2, t0, gp
                                                  30'd    8254    : data = 32'h    00BD3833    ;    //    sltu x16 x26 x11      ====        sltu a6, s10, a1
                                                  30'd    8255    : data = 32'h    01FD8EB3    ;    //    add x29 x27 x31      ====        add t4, s11, t6
                                                  30'd    8256    : data = 32'h    0D1C6713    ;    //    ori x14 x24 209      ====        ori a4, s8, 209
                                                  30'd    8257    : data = 32'h    C71E4313    ;    //    xori x6 x28 -911      ====        xori t1, t3, -911
                                                  30'd    8258    : data = 32'h    015414B3    ;    //    sll x9 x8 x21      ====        sll s1, s0, s5
                                                  30'd    8259    : data = 32'h    63B8CD13    ;    //    xori x26 x17 1595      ====        xori s10, a7, 1595
                                                  30'd    8260    : data = 32'h    01AEA5B3    ;    //    slt x11 x29 x26      ====        slt a1, t4, s10
                                                  30'd    8261    : data = 32'h    014EC9B3    ;    //    xor x19 x29 x20      ====        xor s3, t4, s4
                                                  30'd    8262    : data = 32'h    40930933    ;    //    sub x18 x6 x9      ====        sub s2, t1, s1
                                                  30'd    8263    : data = 32'h    5CD9E8B7    ;    //    lui x17 380318      ====        lui a7, 380318
                                                  30'd    8264    : data = 32'h    A6DA0917    ;    //    auipc x18 683424      ====        auipc s2, 683424
                                                  30'd    8265    : data = 32'h    41545633    ;    //    sra x12 x8 x21      ====        sra a2, s0, s5
                                                  30'd    8266    : data = 32'h    000E05B3    ;    //    add x11 x28 x0      ====        add a1, t3, zero
                                                  30'd    8267    : data = 32'h    61800A97    ;    //    auipc x21 399360      ====        auipc s5, 399360
                                                  30'd    8268    : data = 32'h    4074DB33    ;    //    sra x22 x9 x7      ====        sra s6, s1, t2
                                                  30'd    8269    : data = 32'h    00F6D0B3    ;    //    srl x1 x13 x15      ====        srl ra, a3, a5
                                                  30'd    8270    : data = 32'h    01CFED33    ;    //    or x26 x31 x28      ====        or s10, t6, t3
                                                  30'd    8271    : data = 32'h    01611113    ;    //    slli x2 x2 22      ====        slli sp, sp, 22
                                                  30'd    8272    : data = 32'h    312AAD13    ;    //    slti x26 x21 786      ====        slti s10, s5, 786
                                                  30'd    8273    : data = 32'h    B9442293    ;    //    slti x5 x8 -1132      ====        slti t0, s0, -1132
                                                  30'd    8274    : data = 32'h    40FB5D13    ;    //    srai x26 x22 15      ====        srai s10, s6, 15
                                                  30'd    8275    : data = 32'h    00485E13    ;    //    srli x28 x16 4      ====        srli t3, a6, 4
                                                  30'd    8276    : data = 32'h    EC974313    ;    //    xori x6 x14 -311      ====        xori t1, a4, -311
                                                  30'd    8277    : data = 32'h    21330B93    ;    //    addi x23 x6 531      ====        addi s7, t1, 531
                                                  30'd    8278    : data = 32'h    00A1C8B3    ;    //    xor x17 x3 x10      ====        xor a7, gp, a0
                                                  30'd    8279    : data = 32'h    004FFB33    ;    //    and x22 x31 x4      ====        and s6, t6, tp
                                                  30'd    8280    : data = 32'h    0169CE33    ;    //    xor x28 x19 x22      ====        xor t3, s3, s6
                                                  30'd    8281    : data = 32'h    01984DB3    ;    //    xor x27 x16 x25      ====        xor s11, a6, s9
                                                  30'd    8282    : data = 32'h    0082CBB3    ;    //    xor x23 x5 x8      ====        xor s7, t0, s0
                                                  30'd    8283    : data = 32'h    001B65B3    ;    //    or x11 x22 x1      ====        or a1, s6, ra
                                                  30'd    8284    : data = 32'h    014C3393    ;    //    sltiu x7 x24 20      ====        sltiu t2, s8, 20
                                                  30'd    8285    : data = 32'h    01DDFDB3    ;    //    and x27 x27 x29      ====        and s11, s11, t4
                                                  30'd    8286    : data = 32'h    C37F2B13    ;    //    slti x22 x30 -969      ====        slti s6, t5, -969
                                                  30'd    8287    : data = 32'h    00121D93    ;    //    slli x27 x4 1      ====        slli s11, tp, 1
                                                  30'd    8288    : data = 32'h    00B1BFB3    ;    //    sltu x31 x3 x11      ====        sltu t6, gp, a1
                                                  30'd    8289    : data = 32'h    00C3D2B3    ;    //    srl x5 x7 x12      ====        srl t0, t2, a2
                                                  30'd    8290    : data = 32'h    AD4F3713    ;    //    sltiu x14 x30 -1324      ====        sltiu a4, t5, -1324
                                                  30'd    8291    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8292    : data = 32'h    40E60033    ;    //    sub x0 x12 x14      ====        sub zero, a2, a4
                                                  30'd    8293    : data = 32'h    402086B3    ;    //    sub x13 x1 x2      ====        sub a3, ra, sp
                                                  30'd    8294    : data = 32'h    73420D97    ;    //    auipc x27 472096      ====        auipc s11, 472096
                                                  30'd    8295    : data = 32'h    01A407B3    ;    //    add x15 x8 x26      ====        add a5, s0, s10
                                                  30'd    8296    : data = 32'h    01A9DD33    ;    //    srl x26 x19 x26      ====        srl s10, s3, s10
                                                  30'd    8297    : data = 32'h    01FF70B3    ;    //    and x1 x30 x31      ====        and ra, t5, t6
                                                  30'd    8298    : data = 32'h    E969B393    ;    //    sltiu x7 x19 -362      ====        sltiu t2, s3, -362
                                                  30'd    8299    : data = 32'h    41F956B3    ;    //    sra x13 x18 x31      ====        sra a3, s2, t6
                                                  30'd    8300    : data = 32'h    41A5D893    ;    //    srai x17 x11 26      ====        srai a7, a1, 26
                                                  30'd    8301    : data = 32'h    4140D413    ;    //    srai x8 x1 20      ====        srai s0, ra, 20
                                                  30'd    8302    : data = 32'h    01BDB7B3    ;    //    sltu x15 x27 x27      ====        sltu a5, s11, s11
                                                  30'd    8303    : data = 32'h    40485033    ;    //    sra x0 x16 x4      ====        sra zero, a6, tp
                                                  30'd    8304    : data = 32'h    CBD05717    ;    //    auipc x14 834821      ====        auipc a4, 834821
                                                  30'd    8305    : data = 32'h    9CDD0293    ;    //    addi x5 x26 -1587      ====        addi t0, s10, -1587
                                                  30'd    8306    : data = 32'h    00DC41B3    ;    //    xor x3 x24 x13      ====        xor gp, s8, a3
                                                  30'd    8307    : data = 32'h    AE398137    ;    //    lui x2 713624      ====        lui sp, 713624
                                                  30'd    8308    : data = 32'h    0120D793    ;    //    srli x15 x1 18      ====        srli a5, ra, 18
                                                  30'd    8309    : data = 32'h    01A46633    ;    //    or x12 x8 x26      ====        or a2, s0, s10
                                                  30'd    8310    : data = 32'h    40B783B3    ;    //    sub x7 x15 x11      ====        sub t2, a5, a1
                                                  30'd    8311    : data = 32'h    01A25E33    ;    //    srl x28 x4 x26      ====        srl t3, tp, s10
                                                  30'd    8312    : data = 32'h    B3910B93    ;    //    addi x23 x2 -1223      ====        addi s7, sp, -1223
                                                  30'd    8313    : data = 32'h    EAD5A293    ;    //    slti x5 x11 -339      ====        slti t0, a1, -339
                                                  30'd    8314    : data = 32'h    01C8F333    ;    //    and x6 x17 x28      ====        and t1, a7, t3
                                                  30'd    8315    : data = 32'h    006C0E33    ;    //    add x28 x24 x6      ====        add t3, s8, t1
                                                  30'd    8316    : data = 32'h    6800A493    ;    //    slti x9 x1 1664      ====        slti s1, ra, 1664
                                                  30'd    8317    : data = 32'h    A0A24793    ;    //    xori x15 x4 -1526      ====        xori a5, tp, -1526
                                                  30'd    8318    : data = 32'h    920E6313    ;    //    ori x6 x28 -1760      ====        ori t1, t3, -1760
                                                  30'd    8319    : data = 32'h    E0F5B837    ;    //    lui x16 921435      ====        lui a6, 921435
                                                  30'd    8320    : data = 32'h    487F7613    ;    //    andi x12 x30 1159      ====        andi a2, t5, 1159
                                                  30'd    8321    : data = 32'h    0118DB93    ;    //    srli x23 x17 17      ====        srli s7, a7, 17
                                                  30'd    8322    : data = 32'h    003AFDB3    ;    //    and x27 x21 x3      ====        and s11, s5, gp
                                                  30'd    8323    : data = 32'h    019D0333    ;    //    add x6 x26 x25      ====        add t1, s10, s9
                                                  30'd    8324    : data = 32'h    418600B3    ;    //    sub x1 x12 x24      ====        sub ra, a2, s8
                                                  30'd    8325    : data = 32'h    88614113    ;    //    xori x2 x2 -1914      ====        xori sp, sp, -1914
                                                  30'd    8326    : data = 32'h    41B3D3B3    ;    //    sra x7 x7 x27      ====        sra t2, t2, s11
                                                  30'd    8327    : data = 32'h    01F4AC33    ;    //    slt x24 x9 x31      ====        slt s8, s1, t6
                                                  30'd    8328    : data = 32'h    812AF613    ;    //    andi x12 x21 -2030      ====        andi a2, s5, -2030
                                                  30'd    8329    : data = 32'h    002F11B3    ;    //    sll x3 x30 x2      ====        sll gp, t5, sp
                                                  30'd    8330    : data = 32'h    007709B3    ;    //    add x19 x14 x7      ====        add s3, a4, t2
                                                  30'd    8331    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8332    : data = 32'h    A29DC113    ;    //    xori x2 x27 -1495      ====        xori sp, s11, -1495
                                                  30'd    8333    : data = 32'h    01558D33    ;    //    add x26 x11 x21      ====        add s10, a1, s5
                                                  30'd    8334    : data = 32'h    00CCCBB3    ;    //    xor x23 x25 x12      ====        xor s7, s9, a2
                                                  30'd    8335    : data = 32'h    BEA46293    ;    //    ori x5 x8 -1046      ====        ori t0, s0, -1046
                                                  30'd    8336    : data = 32'h    0069E2B3    ;    //    or x5 x19 x6      ====        or t0, s3, t1
                                                  30'd    8337    : data = 32'h    0129EDB3    ;    //    or x27 x19 x18      ====        or s11, s3, s2
                                                  30'd    8338    : data = 32'h    960C4193    ;    //    xori x3 x24 -1696      ====        xori gp, s8, -1696
                                                  30'd    8339    : data = 32'h    01475EB3    ;    //    srl x29 x14 x20      ====        srl t4, a4, s4
                                                  30'd    8340    : data = 32'h    019F19B3    ;    //    sll x19 x30 x25      ====        sll s3, t5, s9
                                                  30'd    8341    : data = 32'h    00F7C1B3    ;    //    xor x3 x15 x15      ====        xor gp, a5, a5
                                                  30'd    8342    : data = 32'h    01219633    ;    //    sll x12 x3 x18      ====        sll a2, gp, s2
                                                  30'd    8343    : data = 32'h    030EF413    ;    //    andi x8 x29 48      ====        andi s0, t4, 48
                                                  30'd    8344    : data = 32'h    978B6013    ;    //    ori x0 x22 -1672      ====        ori zero, s6, -1672
                                                  30'd    8345    : data = 32'h    009FEB33    ;    //    or x22 x31 x9      ====        or s6, t6, s1
                                                  30'd    8346    : data = 32'h    01FE67B3    ;    //    or x15 x28 x31      ====        or a5, t3, t6
                                                  30'd    8347    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8348    : data = 32'h    01AB23B3    ;    //    slt x7 x22 x26      ====        slt t2, s6, s10
                                                  30'd    8349    : data = 32'h    DD9DB393    ;    //    sltiu x7 x27 -551      ====        sltiu t2, s11, -551
                                                  30'd    8350    : data = 32'h    00D8D733    ;    //    srl x14 x17 x13      ====        srl a4, a7, a3
                                                  30'd    8351    : data = 32'h    00101A13    ;    //    slli x20 x0 1      ====        slli s4, zero, 1
                                                  30'd    8352    : data = 32'h    00BE1D13    ;    //    slli x26 x28 11      ====        slli s10, t3, 11
                                                  30'd    8353    : data = 32'h    AFC7FB13    ;    //    andi x22 x15 -1284      ====        andi s6, a5, -1284
                                                  30'd    8354    : data = 32'h    40670033    ;    //    sub x0 x14 x6      ====        sub zero, a4, t1
                                                  30'd    8355    : data = 32'h    40270A33    ;    //    sub x20 x14 x2      ====        sub s4, a4, sp
                                                  30'd    8356    : data = 32'h    40788133    ;    //    sub x2 x17 x7      ====        sub sp, a7, t2
                                                  30'd    8357    : data = 32'h    40AFD133    ;    //    sra x2 x31 x10      ====        sra sp, t6, a0
                                                  30'd    8358    : data = 32'h    9EC4B793    ;    //    sltiu x15 x9 -1556      ====        sltiu a5, s1, -1556
                                                  30'd    8359    : data = 32'h    014DF733    ;    //    and x14 x27 x20      ====        and a4, s11, s4
                                                  30'd    8360    : data = 32'h    9584AD13    ;    //    slti x26 x9 -1704      ====        slti s10, s1, -1704
                                                  30'd    8361    : data = 32'h    405652B3    ;    //    sra x5 x12 x5      ====        sra t0, a2, t0
                                                  30'd    8362    : data = 32'h    01661013    ;    //    slli x0 x12 22      ====        slli zero, a2, 22
                                                  30'd    8363    : data = 32'h    40460FB3    ;    //    sub x31 x12 x4      ====        sub t6, a2, tp
                                                  30'd    8364    : data = 32'h    00E35793    ;    //    srli x15 x6 14      ====        srli a5, t1, 14
                                                  30'd    8365    : data = 32'h    910EAD13    ;    //    slti x26 x29 -1776      ====        slti s10, t4, -1776
                                                  30'd    8366    : data = 32'h    9AE27D93    ;    //    andi x27 x4 -1618      ====        andi s11, tp, -1618
                                                  30'd    8367    : data = 32'h    33F9B913    ;    //    sltiu x18 x19 831      ====        sltiu s2, s3, 831
                                                  30'd    8368    : data = 32'h    01D55393    ;    //    srli x7 x10 29      ====        srli t2, a0, 29
                                                  30'd    8369    : data = 32'h    E9F8C113    ;    //    xori x2 x17 -353      ====        xori sp, a7, -353
                                                  30'd    8370    : data = 32'h    41BFDFB3    ;    //    sra x31 x31 x27      ====        sra t6, t6, s11
                                                  30'd    8371    : data = 32'h    0166C1B3    ;    //    xor x3 x13 x22      ====        xor gp, a3, s6
                                                  30'd    8372    : data = 32'h    00975EB3    ;    //    srl x29 x14 x9      ====        srl t4, a4, s1
                                                  30'd    8373    : data = 32'h    5ECD3C37    ;    //    lui x24 388307      ====        lui s8, 388307
                                                  30'd    8374    : data = 32'h    ADC7C193    ;    //    xori x3 x15 -1316      ====        xori gp, a5, -1316
                                                  30'd    8375    : data = 32'h    403F8033    ;    //    sub x0 x31 x3      ====        sub zero, t6, gp
                                                  30'd    8376    : data = 32'h    F520D4B7    ;    //    lui x9 1004045      ====        lui s1, 1004045
                                                  30'd    8377    : data = 32'h    ED88E793    ;    //    ori x15 x17 -296      ====        ori a5, a7, -296
                                                  30'd    8378    : data = 32'h    01F562B3    ;    //    or x5 x10 x31      ====        or t0, a0, t6
                                                  30'd    8379    : data = 32'h    40EB5813    ;    //    srai x16 x22 14      ====        srai a6, s6, 14
                                                  30'd    8380    : data = 32'h    C1BC4613    ;    //    xori x12 x24 -997      ====        xori a2, s8, -997
                                                  30'd    8381    : data = 32'h    6DBCEC93    ;    //    ori x25 x25 1755      ====        ori s9, s9, 1755
                                                  30'd    8382    : data = 32'h    00734733    ;    //    xor x14 x6 x7      ====        xor a4, t1, t2
                                                  30'd    8383    : data = 32'h    41628433    ;    //    sub x8 x5 x22      ====        sub s0, t0, s6
                                                  30'd    8384    : data = 32'h    00B95633    ;    //    srl x12 x18 x11      ====        srl a2, s2, a1
                                                  30'd    8385    : data = 32'h    B0A20F93    ;    //    addi x31 x4 -1270      ====        addi t6, tp, -1270
                                                  30'd    8386    : data = 32'h    00D02D33    ;    //    slt x26 x0 x13      ====        slt s10, zero, a3
                                                  30'd    8387    : data = 32'h    0051CB33    ;    //    xor x22 x3 x5      ====        xor s6, gp, t0
                                                  30'd    8388    : data = 32'h    41D05A13    ;    //    srai x20 x0 29      ====        srai s4, zero, 29
                                                  30'd    8389    : data = 32'h    D3D22413    ;    //    slti x8 x4 -707      ====        slti s0, tp, -707
                                                  30'd    8390    : data = 32'h    00DD46B3    ;    //    xor x13 x26 x13      ====        xor a3, s10, a3
                                                  30'd    8391    : data = 32'h    012524B3    ;    //    slt x9 x10 x18      ====        slt s1, a0, s2
                                                  30'd    8392    : data = 32'h    41B05493    ;    //    srai x9 x0 27      ====        srai s1, zero, 27
                                                  30'd    8393    : data = 32'h    41AFD413    ;    //    srai x8 x31 26      ====        srai s0, t6, 26
                                                  30'd    8394    : data = 32'h    954A7193    ;    //    andi x3 x20 -1708      ====        andi gp, s4, -1708
                                                  30'd    8395    : data = 32'h    00814433    ;    //    xor x8 x2 x8      ====        xor s0, sp, s0
                                                  30'd    8396    : data = 32'h    254E4813    ;    //    xori x16 x28 596      ====        xori a6, t3, 596
                                                  30'd    8397    : data = 32'h    01936A33    ;    //    or x20 x6 x25      ====        or s4, t1, s9
                                                  30'd    8398    : data = 32'h    018F6033    ;    //    or x0 x30 x24      ====        or zero, t5, s8
                                                  30'd    8399    : data = 32'h    C4CA4117    ;    //    auipc x2 806052      ====        auipc sp, 806052
                                                  30'd    8400    : data = 32'h    00F5DD93    ;    //    srli x27 x11 15      ====        srli s11, a1, 15
                                                  30'd    8401    : data = 32'h    8CE5E337    ;    //    lui x6 577118      ====        lui t1, 577118
                                                  30'd    8402    : data = 32'h    00BF60B3    ;    //    or x1 x30 x11      ====        or ra, t5, a1
                                                  30'd    8403    : data = 32'h    22604713    ;    //    xori x14 x0 550      ====        xori a4, zero, 550
                                                  30'd    8404    : data = 32'h    99EA4A13    ;    //    xori x20 x20 -1634      ====        xori s4, s4, -1634
                                                  30'd    8405    : data = 32'h    405A0BB3    ;    //    sub x23 x20 x5      ====        sub s7, s4, t0
                                                  30'd    8406    : data = 32'h    C2E794B7    ;    //    lui x9 798329      ====        lui s1, 798329
                                                  30'd    8407    : data = 32'h    7B6CBB13    ;    //    sltiu x22 x25 1974      ====        sltiu s6, s9, 1974
                                                  30'd    8408    : data = 32'h    01F17B33    ;    //    and x22 x2 x31      ====        and s6, sp, t6
                                                  30'd    8409    : data = 32'h    00E3A2B3    ;    //    slt x5 x7 x14      ====        slt t0, t2, a4
                                                  30'd    8410    : data = 32'h    CC0E3093    ;    //    sltiu x1 x28 -832      ====        sltiu ra, t3, -832
                                                  30'd    8411    : data = 32'h    01CE7FB3    ;    //    and x31 x28 x28      ====        and t6, t3, t3
                                                  30'd    8412    : data = 32'h    003A42B3    ;    //    xor x5 x20 x3      ====        xor t0, s4, gp
                                                  30'd    8413    : data = 32'h    01A03D33    ;    //    sltu x26 x0 x26      ====        sltu s10, zero, s10
                                                  30'd    8414    : data = 32'h    6454D797    ;    //    auipc x15 410957      ====        auipc a5, 410957
                                                  30'd    8415    : data = 32'h    0F2CC593    ;    //    xori x11 x25 242      ====        xori a1, s9, 242
                                                  30'd    8416    : data = 32'h    418DD313    ;    //    srai x6 x27 24      ====        srai t1, s11, 24
                                                  30'd    8417    : data = 32'h    21C5C6B7    ;    //    lui x13 138332      ====        lui a3, 138332
                                                  30'd    8418    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8419    : data = 32'h    410ADB13    ;    //    srai x22 x21 16      ====        srai s6, s5, 16
                                                  30'd    8420    : data = 32'h    004D5813    ;    //    srli x16 x26 4      ====        srli a6, s10, 4
                                                  30'd    8421    : data = 32'h    41078A33    ;    //    sub x20 x15 x16      ====        sub s4, a5, a6
                                                  30'd    8422    : data = 32'h    002670B3    ;    //    and x1 x12 x2      ====        and ra, a2, sp
                                                  30'd    8423    : data = 32'h    EBB24A13    ;    //    xori x20 x4 -325      ====        xori s4, tp, -325
                                                  30'd    8424    : data = 32'h    00C99CB3    ;    //    sll x25 x19 x12      ====        sll s9, s3, a2
                                                  30'd    8425    : data = 32'h    00C0DE93    ;    //    srli x29 x1 12      ====        srli t4, ra, 12
                                                  30'd    8426    : data = 32'h    00DA5D13    ;    //    srli x26 x20 13      ====        srli s10, s4, 13
                                                  30'd    8427    : data = 32'h    01031633    ;    //    sll x12 x6 x16      ====        sll a2, t1, a6
                                                  30'd    8428    : data = 32'h    41D80033    ;    //    sub x0 x16 x29      ====        sub zero, a6, t4
                                                  30'd    8429    : data = 32'h    2096B793    ;    //    sltiu x15 x13 521      ====        sltiu a5, a3, 521
                                                  30'd    8430    : data = 32'h    01731493    ;    //    slli x9 x6 23      ====        slli s1, t1, 23
                                                  30'd    8431    : data = 32'h    000CDE93    ;    //    srli x29 x25 0      ====        srli t4, s9, 0
                                                  30'd    8432    : data = 32'h    A3632137    ;    //    lui x2 669234      ====        lui sp, 669234
                                                  30'd    8433    : data = 32'h    40C75693    ;    //    srai x13 x14 12      ====        srai a3, a4, 12
                                                  30'd    8434    : data = 32'h    4B5A8F93    ;    //    addi x31 x21 1205      ====        addi t6, s5, 1205
                                                  30'd    8435    : data = 32'h    75DCBB17    ;    //    auipc x22 482763      ====        auipc s6, 482763
                                                  30'd    8436    : data = 32'h    00154EB3    ;    //    xor x29 x10 x1      ====        xor t4, a0, ra
                                                  30'd    8437    : data = 32'h    4106DEB3    ;    //    sra x29 x13 x16      ====        sra t4, a3, a6
                                                  30'd    8438    : data = 32'h    013286B3    ;    //    add x13 x5 x19      ====        add a3, t0, s3
                                                  30'd    8439    : data = 32'h    5D97E917    ;    //    auipc x18 383358      ====        auipc s2, 383358
                                                  30'd    8440    : data = 32'h    83BA7C13    ;    //    andi x24 x20 -1989      ====        andi s8, s4, -1989
                                                  30'd    8441    : data = 32'h    2FDC0637    ;    //    lui x12 196032      ====        lui a2, 196032
                                                  30'd    8442    : data = 32'h    41B5DA33    ;    //    sra x20 x11 x27      ====        sra s4, a1, s11
                                                  30'd    8443    : data = 32'h    01DB0EB3    ;    //    add x29 x22 x29      ====        add t4, s6, t4
                                                  30'd    8444    : data = 32'h    B4B93613    ;    //    sltiu x12 x18 -1205      ====        sltiu a2, s2, -1205
                                                  30'd    8445    : data = 32'h    00F776B3    ;    //    and x13 x14 x15      ====        and a3, a4, a5
                                                  30'd    8446    : data = 32'h    D0BD4B13    ;    //    xori x22 x26 -757      ====        xori s6, s10, -757
                                                  30'd    8447    : data = 32'h    EEC42D13    ;    //    slti x26 x8 -276      ====        slti s10, s0, -276
                                                  30'd    8448    : data = 32'h    41E482B3    ;    //    sub x5 x9 x30      ====        sub t0, s1, t5
                                                  30'd    8449    : data = 32'h    40F25C93    ;    //    srai x25 x4 15      ====        srai s9, tp, 15
                                                  30'd    8450    : data = 32'h    41D15A13    ;    //    srai x20 x2 29      ====        srai s4, sp, 29
                                                  30'd    8451    : data = 32'h    401981B3    ;    //    sub x3 x19 x1      ====        sub gp, s3, ra
                                                  30'd    8452    : data = 32'h    013BB7B3    ;    //    sltu x15 x23 x19      ====        sltu a5, s7, s3
                                                  30'd    8453    : data = 32'h    00310B33    ;    //    add x22 x2 x3      ====        add s6, sp, gp
                                                  30'd    8454    : data = 32'h    0124BE33    ;    //    sltu x28 x9 x18      ====        sltu t3, s1, s2
                                                  30'd    8455    : data = 32'h    FB27A313    ;    //    slti x6 x15 -78      ====        slti t1, a5, -78
                                                  30'd    8456    : data = 32'h    0089BDB3    ;    //    sltu x27 x19 x8      ====        sltu s11, s3, s0
                                                  30'd    8457    : data = 32'h    3A83F293    ;    //    andi x5 x7 936      ====        andi t0, t2, 936
                                                  30'd    8458    : data = 32'h    00635193    ;    //    srli x3 x6 6      ====        srli gp, t1, 6
                                                  30'd    8459    : data = 32'h    01C6D033    ;    //    srl x0 x13 x28      ====        srl zero, a3, t3
                                                  30'd    8460    : data = 32'h    AE4FB893    ;    //    sltiu x17 x31 -1308      ====        sltiu a7, t6, -1308
                                                  30'd    8461    : data = 32'h    026FC913    ;    //    xori x18 x31 38      ====        xori s2, t6, 38
                                                  30'd    8462    : data = 32'h    01B27D33    ;    //    and x26 x4 x27      ====        and s10, tp, s11
                                                  30'd    8463    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8464    : data = 32'h    4163D913    ;    //    srai x18 x7 22      ====        srai s2, t2, 22
                                                  30'd    8465    : data = 32'h    009B2433    ;    //    slt x8 x22 x9      ====        slt s0, s6, s1
                                                  30'd    8466    : data = 32'h    01B53633    ;    //    sltu x12 x10 x27      ====        sltu a2, a0, s11
                                                  30'd    8467    : data = 32'h    F63C4C13    ;    //    xori x24 x24 -157      ====        xori s8, s8, -157
                                                  30'd    8468    : data = 32'h    40345C13    ;    //    srai x24 x8 3      ====        srai s8, s0, 3
                                                  30'd    8469    : data = 32'h    0D554113    ;    //    xori x2 x10 213      ====        xori sp, a0, 213
                                                  30'd    8470    : data = 32'h    01FAB333    ;    //    sltu x6 x21 x31      ====        sltu t1, s5, t6
                                                  30'd    8471    : data = 32'h    469B0293    ;    //    addi x5 x22 1129      ====        addi t0, s6, 1129
                                                  30'd    8472    : data = 32'h    01CC61B3    ;    //    or x3 x24 x28      ====        or gp, s8, t3
                                                  30'd    8473    : data = 32'h    BF0D7613    ;    //    andi x12 x26 -1040      ====        andi a2, s10, -1040
                                                  30'd    8474    : data = 32'h    0014E333    ;    //    or x6 x9 x1      ====        or t1, s1, ra
                                                  30'd    8475    : data = 32'h    241D9117    ;    //    auipc x2 147929      ====        auipc sp, 147929
                                                  30'd    8476    : data = 32'h    002D9833    ;    //    sll x16 x27 x2      ====        sll a6, s11, sp
                                                  30'd    8477    : data = 32'h    45BBC097    ;    //    auipc x1 285628      ====        auipc ra, 285628
                                                  30'd    8478    : data = 32'h    009B2433    ;    //    slt x8 x22 x9      ====        slt s0, s6, s1
                                                  30'd    8479    : data = 32'h    77E70093    ;    //    addi x1 x14 1918      ====        addi ra, a4, 1918
                                                  30'd    8480    : data = 32'h    00C2F5B3    ;    //    and x11 x5 x12      ====        and a1, t0, a2
                                                  30'd    8481    : data = 32'h    011C0DB3    ;    //    add x27 x24 x17      ====        add s11, s8, a7
                                                  30'd    8482    : data = 32'h    01202DB3    ;    //    slt x27 x0 x18      ====        slt s11, zero, s2
                                                  30'd    8483    : data = 32'h    40638933    ;    //    sub x18 x7 x6      ====        sub s2, t2, t1
                                                  30'd    8484    : data = 32'h    D8F67E13    ;    //    andi x28 x12 -625      ====        andi t3, a2, -625
                                                  30'd    8485    : data = 32'h    C4B6B913    ;    //    sltiu x18 x13 -949      ====        sltiu s2, a3, -949
                                                  30'd    8486    : data = 32'h    58337D13    ;    //    andi x26 x6 1411      ====        andi s10, t1, 1411
                                                  30'd    8487    : data = 32'h    00D158B3    ;    //    srl x17 x2 x13      ====        srl a7, sp, a3
                                                  30'd    8488    : data = 32'h    26CBBB13    ;    //    sltiu x22 x23 620      ====        sltiu s6, s7, 620
                                                  30'd    8489    : data = 32'h    0123C4B3    ;    //    xor x9 x7 x18      ====        xor s1, t2, s2
                                                  30'd    8490    : data = 32'h    BF2C0DB7    ;    //    lui x27 783040      ====        lui s11, 783040
                                                  30'd    8491    : data = 32'h    40558C33    ;    //    sub x24 x11 x5      ====        sub s8, a1, t0
                                                  30'd    8492    : data = 32'h    8A120893    ;    //    addi x17 x4 -1887      ====        addi a7, tp, -1887
                                                  30'd    8493    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8494    : data = 32'h    41600B33    ;    //    sub x22 x0 x22      ====        sub s6, zero, s6
                                                  30'd    8495    : data = 32'h    01E8A033    ;    //    slt x0 x17 x30      ====        slt zero, a7, t5
                                                  30'd    8496    : data = 32'h    00714FB3    ;    //    xor x31 x2 x7      ====        xor t6, sp, t2
                                                  30'd    8497    : data = 32'h    00E78AB3    ;    //    add x21 x15 x14      ====        add s5, a5, a4
                                                  30'd    8498    : data = 32'h    0190CDB3    ;    //    xor x27 x1 x25      ====        xor s11, ra, s9
                                                  30'd    8499    : data = 32'h    D82C4893    ;    //    xori x17 x24 -638      ====        xori a7, s8, -638
                                                  30'd    8500    : data = 32'h    406BD6B3    ;    //    sra x13 x23 x6      ====        sra a3, s7, t1
                                                  30'd    8501    : data = 32'h    B0D4DA97    ;    //    auipc x21 724301      ====        auipc s5, 724301
                                                  30'd    8502    : data = 32'h    63D7D417    ;    //    auipc x8 408957      ====        auipc s0, 408957
                                                  30'd    8503    : data = 32'h    01704AB3    ;    //    xor x21 x0 x23      ====        xor s5, zero, s7
                                                  30'd    8504    : data = 32'h    4058D033    ;    //    sra x0 x17 x5      ====        sra zero, a7, t0
                                                  30'd    8505    : data = 32'h    000D1FB3    ;    //    sll x31 x26 x0      ====        sll t6, s10, zero
                                                  30'd    8506    : data = 32'h    DD5D62B7    ;    //    lui x5 906710      ====        lui t0, 906710
                                                  30'd    8507    : data = 32'h    40AA5713    ;    //    srai x14 x20 10      ====        srai a4, s4, 10
                                                  30'd    8508    : data = 32'h    01E5DE93    ;    //    srli x29 x11 30      ====        srli t4, a1, 30
                                                  30'd    8509    : data = 32'h    89810413    ;    //    addi x8 x2 -1896      ====        addi s0, sp, -1896
                                                  30'd    8510    : data = 32'h    4146D0B3    ;    //    sra x1 x13 x20      ====        sra ra, a3, s4
                                                  30'd    8511    : data = 32'h    01B033B3    ;    //    sltu x7 x0 x27      ====        sltu t2, zero, s11
                                                  30'd    8512    : data = 32'h    48640913    ;    //    addi x18 x8 1158      ====        addi s2, s0, 1158
                                                  30'd    8513    : data = 32'h    36104913    ;    //    xori x18 x0 865      ====        xori s2, zero, 865
                                                  30'd    8514    : data = 32'h    01FDCD33    ;    //    xor x26 x27 x31      ====        xor s10, s11, t6
                                                  30'd    8515    : data = 32'h    F5897C93    ;    //    andi x25 x18 -168      ====        andi s9, s2, -168
                                                  30'd    8516    : data = 32'h    00D3A2B3    ;    //    slt x5 x7 x13      ====        slt t0, t2, a3
                                                  30'd    8517    : data = 32'h    01785413    ;    //    srli x8 x16 23      ====        srli s0, a6, 23
                                                  30'd    8518    : data = 32'h    0174BB33    ;    //    sltu x22 x9 x23      ====        sltu s6, s1, s7
                                                  30'd    8519    : data = 32'h    00EE9E93    ;    //    slli x29 x29 14      ====        slli t4, t4, 14
                                                  30'd    8520    : data = 32'h    DFDBFC17    ;    //    auipc x24 916927      ====        auipc s8, 916927
                                                  30'd    8521    : data = 32'h    40355293    ;    //    srai x5 x10 3      ====        srai t0, a0, 3
                                                  30'd    8522    : data = 32'h    CEF0EB97    ;    //    auipc x23 847630      ====        auipc s7, 847630
                                                  30'd    8523    : data = 32'h    00CA1D13    ;    //    slli x26 x20 12      ====        slli s10, s4, 12
                                                  30'd    8524    : data = 32'h    004E1293    ;    //    slli x5 x28 4      ====        slli t0, t3, 4
                                                  30'd    8525    : data = 32'h    00259B93    ;    //    slli x23 x11 2      ====        slli s7, a1, 2
                                                  30'd    8526    : data = 32'h    0CC37A13    ;    //    andi x20 x6 204      ====        andi s4, t1, 204
                                                  30'd    8527    : data = 32'h    41725893    ;    //    srai x17 x4 23      ====        srai a7, tp, 23
                                                  30'd    8528    : data = 32'h    00DB1C93    ;    //    slli x25 x22 13      ====        slli s9, s6, 13
                                                  30'd    8529    : data = 32'h    00CAB4B3    ;    //    sltu x9 x21 x12      ====        sltu s1, s5, a2
                                                  30'd    8530    : data = 32'h    4025DE33    ;    //    sra x28 x11 x2      ====        sra t3, a1, sp
                                                  30'd    8531    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8532    : data = 32'h    00E478B3    ;    //    and x17 x8 x14      ====        and a7, s0, a4
                                                  30'd    8533    : data = 32'h    40C281B3    ;    //    sub x3 x5 x12      ====        sub gp, t0, a2
                                                  30'd    8534    : data = 32'h    0075EE33    ;    //    or x28 x11 x7      ====        or t3, a1, t2
                                                  30'd    8535    : data = 32'h    01831793    ;    //    slli x15 x6 24      ====        slli a5, t1, 24
                                                  30'd    8536    : data = 32'h    FFEEF393    ;    //    andi x7 x29 -2      ====        andi t2, t4, -2
                                                  30'd    8537    : data = 32'h    019D9E33    ;    //    sll x28 x27 x25      ====        sll t3, s11, s9
                                                  30'd    8538    : data = 32'h    0164CC33    ;    //    xor x24 x9 x22      ====        xor s8, s1, s6
                                                  30'd    8539    : data = 32'h    0162C0B3    ;    //    xor x1 x5 x22      ====        xor ra, t0, s6
                                                  30'd    8540    : data = 32'h    2E6BA393    ;    //    slti x7 x23 742      ====        slti t2, s7, 742
                                                  30'd    8541    : data = 32'h    003391B3    ;    //    sll x3 x7 x3      ====        sll gp, t2, gp
                                                  30'd    8542    : data = 32'h    407E0AB3    ;    //    sub x21 x28 x7      ====        sub s5, t3, t2
                                                  30'd    8543    : data = 32'h    01BD2033    ;    //    slt x0 x26 x27      ====        slt zero, s10, s11
                                                  30'd    8544    : data = 32'h    9E492C17    ;    //    auipc x24 648338      ====        auipc s8, 648338
                                                  30'd    8545    : data = 32'h    B5330293    ;    //    addi x5 x6 -1197      ====        addi t0, t1, -1197
                                                  30'd    8546    : data = 32'h    41F002B3    ;    //    sub x5 x0 x31      ====        sub t0, zero, t6
                                                  30'd    8547    : data = 32'h    6C0684B7    ;    //    lui x9 442472      ====        lui s1, 442472
                                                  30'd    8548    : data = 32'h    926A4C13    ;    //    xori x24 x20 -1754      ====        xori s8, s4, -1754
                                                  30'd    8549    : data = 32'h    01E45393    ;    //    srli x7 x8 30      ====        srli t2, s0, 30
                                                  30'd    8550    : data = 32'h    0006E7B3    ;    //    or x15 x13 x0      ====        or a5, a3, zero
                                                  30'd    8551    : data = 32'h    2F09AA93    ;    //    slti x21 x19 752      ====        slti s5, s3, 752
                                                  30'd    8552    : data = 32'h    FF8B38B7    ;    //    lui x17 1046707      ====        lui a7, 1046707
                                                  30'd    8553    : data = 32'h    4066D033    ;    //    sra x0 x13 x6      ====        sra zero, a3, t1
                                                  30'd    8554    : data = 32'h    007EEBB3    ;    //    or x23 x29 x7      ====        or s7, t4, t2
                                                  30'd    8555    : data = 32'h    6FF34F97    ;    //    auipc x31 458548      ====        auipc t6, 458548
                                                  30'd    8556    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8557    : data = 32'h    01847733    ;    //    and x14 x8 x24      ====        and a4, s0, s8
                                                  30'd    8558    : data = 32'h    41DF5313    ;    //    srai x6 x30 29      ====        srai t1, t5, 29
                                                  30'd    8559    : data = 32'h    00B68133    ;    //    add x2 x13 x11      ====        add sp, a3, a1
                                                  30'd    8560    : data = 32'h    C4982793    ;    //    slti x15 x16 -951      ====        slti a5, a6, -951
                                                  30'd    8561    : data = 32'h    000CCE33    ;    //    xor x28 x25 x0      ====        xor t3, s9, zero
                                                  30'd    8562    : data = 32'h    60D06093    ;    //    ori x1 x0 1549      ====        ori ra, zero, 1549
                                                  30'd    8563    : data = 32'h    39DC4313    ;    //    xori x6 x24 925      ====        xori t1, s8, 925
                                                  30'd    8564    : data = 32'h    E8141437    ;    //    lui x8 950593      ====        lui s0, 950593
                                                  30'd    8565    : data = 32'h    01A7B333    ;    //    sltu x6 x15 x26      ====        sltu t1, a5, s10
                                                  30'd    8566    : data = 32'h    012E9933    ;    //    sll x18 x29 x18      ====        sll s2, t4, s2
                                                  30'd    8567    : data = 32'h    018DD133    ;    //    srl x2 x27 x24      ====        srl sp, s11, s8
                                                  30'd    8568    : data = 32'h    018AC5B3    ;    //    xor x11 x21 x24      ====        xor a1, s5, s8
                                                  30'd    8569    : data = 32'h    0CA9D917    ;    //    auipc x18 51869      ====        auipc s2, 51869
                                                  30'd    8570    : data = 32'h    00E3C2B3    ;    //    xor x5 x7 x14      ====        xor t0, t2, a4
                                                  30'd    8571    : data = 32'h    00B80E33    ;    //    add x28 x16 x11      ====        add t3, a6, a1
                                                  30'd    8572    : data = 32'h    41BDDA13    ;    //    srai x20 x27 27      ====        srai s4, s11, 27
                                                  30'd    8573    : data = 32'h    FB023997    ;    //    auipc x19 1028131      ====        auipc s3, 1028131
                                                  30'd    8574    : data = 32'h    6290E793    ;    //    ori x15 x1 1577      ====        ori a5, ra, 1577
                                                  30'd    8575    : data = 32'h    40B3D433    ;    //    sra x8 x7 x11      ====        sra s0, t2, a1
                                                  30'd    8576    : data = 32'h    7112CD13    ;    //    xori x26 x5 1809      ====        xori s10, t0, 1809
                                                  30'd    8577    : data = 32'h    010668B3    ;    //    or x17 x12 x16      ====        or a7, a2, a6
                                                  30'd    8578    : data = 32'h    58CEAC93    ;    //    slti x25 x29 1420      ====        slti s9, t4, 1420
                                                  30'd    8579    : data = 32'h    017E6133    ;    //    or x2 x28 x23      ====        or sp, t3, s7
                                                  30'd    8580    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8581    : data = 32'h    41CE5413    ;    //    srai x8 x28 28      ====        srai s0, t3, 28
                                                  30'd    8582    : data = 32'h    C95C8D13    ;    //    addi x26 x25 -875      ====        addi s10, s9, -875
                                                  30'd    8583    : data = 32'h    01EF0833    ;    //    add x16 x30 x30      ====        add a6, t5, t5
                                                  30'd    8584    : data = 32'h    00D02E33    ;    //    slt x28 x0 x13      ====        slt t3, zero, a3
                                                  30'd    8585    : data = 32'h    40950133    ;    //    sub x2 x10 x9      ====        sub sp, a0, s1
                                                  30'd    8586    : data = 32'h    00972933    ;    //    slt x18 x14 x9      ====        slt s2, a4, s1
                                                  30'd    8587    : data = 32'h    000A5E13    ;    //    srli x28 x20 0      ====        srli t3, s4, 0
                                                  30'd    8588    : data = 32'h    40FED193    ;    //    srai x3 x29 15      ====        srai gp, t4, 15
                                                  30'd    8589    : data = 32'h    003F5113    ;    //    srli x2 x30 3      ====        srli sp, t5, 3
                                                  30'd    8590    : data = 32'h    005C63B3    ;    //    or x7 x24 x5      ====        or t2, s8, t0
                                                  30'd    8591    : data = 32'h    01C23E33    ;    //    sltu x28 x4 x28      ====        sltu t3, tp, t3
                                                  30'd    8592    : data = 32'h    8FD07A13    ;    //    andi x20 x0 -1795      ====        andi s4, zero, -1795
                                                  30'd    8593    : data = 32'h    E1298C93    ;    //    addi x25 x19 -494      ====        addi s9, s3, -494
                                                  30'd    8594    : data = 32'h    1AF9E817    ;    //    auipc x16 110494      ====        auipc a6, 110494
                                                  30'd    8595    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8596    : data = 32'h    05C80D93    ;    //    addi x27 x16 92      ====        addi s11, a6, 92
                                                  30'd    8597    : data = 32'h    004ACAB3    ;    //    xor x21 x21 x4      ====        xor s5, s5, tp
                                                  30'd    8598    : data = 32'h    00339B93    ;    //    slli x23 x7 3      ====        slli s7, t2, 3
                                                  30'd    8599    : data = 32'h    011D5133    ;    //    srl x2 x26 x17      ====        srl sp, s10, a7
                                                  30'd    8600    : data = 32'h    001508B3    ;    //    add x17 x10 x1      ====        add a7, a0, ra
                                                  30'd    8601    : data = 32'h    41B28EB3    ;    //    sub x29 x5 x27      ====        sub t4, t0, s11
                                                  30'd    8602    : data = 32'h    00E9A0B3    ;    //    slt x1 x19 x14      ====        slt ra, s3, a4
                                                  30'd    8603    : data = 32'h    00B75413    ;    //    srli x8 x14 11      ====        srli s0, a4, 11
                                                  30'd    8604    : data = 32'h    008F58B3    ;    //    srl x17 x30 x8      ====        srl a7, t5, s0
                                                  30'd    8605    : data = 32'h    000F90B3    ;    //    sll x1 x31 x0      ====        sll ra, t6, zero
                                                  30'd    8606    : data = 32'h    01A89493    ;    //    slli x9 x17 26      ====        slli s1, a7, 26
                                                  30'd    8607    : data = 32'h    416A0E33    ;    //    sub x28 x20 x22      ====        sub t3, s4, s6
                                                  30'd    8608    : data = 32'h    00397433    ;    //    and x8 x18 x3      ====        and s0, s2, gp
                                                  30'd    8609    : data = 32'h    00ECD193    ;    //    srli x3 x25 14      ====        srli gp, s9, 14
                                                  30'd    8610    : data = 32'h    3567F013    ;    //    andi x0 x15 854      ====        andi zero, a5, 854
                                                  30'd    8611    : data = 32'h    017D9D13    ;    //    slli x26 x27 23      ====        slli s10, s11, 23
                                                  30'd    8612    : data = 32'h    00A46A33    ;    //    or x20 x8 x10      ====        or s4, s0, a0
                                                  30'd    8613    : data = 32'h    021A3B37    ;    //    lui x22 8611      ====        lui s6, 8611
                                                  30'd    8614    : data = 32'h    01121B93    ;    //    slli x23 x4 17      ====        slli s7, tp, 17
                                                  30'd    8615    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8616    : data = 32'h    C2EA6F93    ;    //    ori x31 x20 -978      ====        ori t6, s4, -978
                                                  30'd    8617    : data = 32'h    D4CE6C93    ;    //    ori x25 x28 -692      ====        ori s9, t3, -692
                                                  30'd    8618    : data = 32'h    B1796937    ;    //    lui x18 726934      ====        lui s2, 726934
                                                  30'd    8619    : data = 32'h    B5720793    ;    //    addi x15 x4 -1193      ====        addi a5, tp, -1193
                                                  30'd    8620    : data = 32'h    097FC713    ;    //    xori x14 x31 151      ====        xori a4, t6, 151
                                                  30'd    8621    : data = 32'h    419106B3    ;    //    sub x13 x2 x25      ====        sub a3, sp, s9
                                                  30'd    8622    : data = 32'h    012D6633    ;    //    or x12 x26 x18      ====        or a2, s10, s2
                                                  30'd    8623    : data = 32'h    6D20AA37    ;    //    lui x20 446986      ====        lui s4, 446986
                                                  30'd    8624    : data = 32'h    04792913    ;    //    slti x18 x18 71      ====        slti s2, s2, 71
                                                  30'd    8625    : data = 32'h    0038C033    ;    //    xor x0 x17 x3      ====        xor zero, a7, gp
                                                  30'd    8626    : data = 32'h    0A1A6197    ;    //    auipc x3 41382      ====        auipc gp, 41382
                                                  30'd    8627    : data = 32'h    01665433    ;    //    srl x8 x12 x22      ====        srl s0, a2, s6
                                                  30'd    8628    : data = 32'h    2F503C93    ;    //    sltiu x25 x0 757      ====        sltiu s9, zero, 757
                                                  30'd    8629    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8630    : data = 32'h    1A0D7E13    ;    //    andi x28 x26 416      ====        andi t3, s10, 416
                                                  30'd    8631    : data = 32'h    001CDB33    ;    //    srl x22 x25 x1      ====        srl s6, s9, ra
                                                  30'd    8632    : data = 32'h    55E48337    ;    //    lui x6 351816      ====        lui t1, 351816
                                                  30'd    8633    : data = 32'h    9D077193    ;    //    andi x3 x14 -1584      ====        andi gp, a4, -1584
                                                  30'd    8634    : data = 32'h    01A82833    ;    //    slt x16 x16 x26      ====        slt a6, a6, s10
                                                  30'd    8635    : data = 32'h    62C1CA93    ;    //    xori x21 x3 1580      ====        xori s5, gp, 1580
                                                  30'd    8636    : data = 32'h    007AF633    ;    //    and x12 x21 x7      ====        and a2, s5, t2
                                                  30'd    8637    : data = 32'h    D35BCD17    ;    //    auipc x26 865724      ====        auipc s10, 865724
                                                  30'd    8638    : data = 32'h    00A99733    ;    //    sll x14 x19 x10      ====        sll a4, s3, a0
                                                  30'd    8639    : data = 32'h    01C7FC33    ;    //    and x24 x15 x28      ====        and s8, a5, t3
                                                  30'd    8640    : data = 32'h    41528733    ;    //    sub x14 x5 x21      ====        sub a4, t0, s5
                                                  30'd    8641    : data = 32'h    BB5F4813    ;    //    xori x16 x30 -1099      ====        xori a6, t5, -1099
                                                  30'd    8642    : data = 32'h    764A6F97    ;    //    auipc x31 484518      ====        auipc t6, 484518
                                                  30'd    8643    : data = 32'h    40E0D393    ;    //    srai x7 x1 14      ====        srai t2, ra, 14
                                                  30'd    8644    : data = 32'h    01D09AB3    ;    //    sll x21 x1 x29      ====        sll s5, ra, t4
                                                  30'd    8645    : data = 32'h    01037D33    ;    //    and x26 x6 x16      ====        and s10, t1, a6
                                                  30'd    8646    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8647    : data = 32'h    00CA9293    ;    //    slli x5 x21 12      ====        slli t0, s5, 12
                                                  30'd    8648    : data = 32'h    014F5E33    ;    //    srl x28 x30 x20      ====        srl t3, t5, s4
                                                  30'd    8649    : data = 32'h    ABE7C413    ;    //    xori x8 x15 -1346      ====        xori s0, a5, -1346
                                                  30'd    8650    : data = 32'h    0106DC13    ;    //    srli x24 x13 16      ====        srli s8, a3, 16
                                                  30'd    8651    : data = 32'h    010276B3    ;    //    and x13 x4 x16      ====        and a3, tp, a6
                                                  30'd    8652    : data = 32'h    00F19D33    ;    //    sll x26 x3 x15      ====        sll s10, gp, a5
                                                  30'd    8653    : data = 32'h    40DBD433    ;    //    sra x8 x23 x13      ====        sra s0, s7, a3
                                                  30'd    8654    : data = 32'h    E0FE0793    ;    //    addi x15 x28 -497      ====        addi a5, t3, -497
                                                  30'd    8655    : data = 32'h    89EE6593    ;    //    ori x11 x28 -1890      ====        ori a1, t3, -1890
                                                  30'd    8656    : data = 32'h    F9064193    ;    //    xori x3 x12 -112      ====        xori gp, a2, -112
                                                  30'd    8657    : data = 32'h    0101A333    ;    //    slt x6 x3 x16      ====        slt t1, gp, a6
                                                  30'd    8658    : data = 32'h    72083713    ;    //    sltiu x14 x16 1824      ====        sltiu a4, a6, 1824
                                                  30'd    8659    : data = 32'h    418FD4B3    ;    //    sra x9 x31 x24      ====        sra s1, t6, s8
                                                  30'd    8660    : data = 32'h    40BF02B3    ;    //    sub x5 x30 x11      ====        sub t0, t5, a1
                                                  30'd    8661    : data = 32'h    D439B9B7    ;    //    lui x19 869275      ====        lui s3, 869275
                                                  30'd    8662    : data = 32'h    51E7AE13    ;    //    slti x28 x15 1310      ====        slti t3, a5, 1310
                                                  30'd    8663    : data = 32'h    ADAADAB7    ;    //    lui x21 711341      ====        lui s5, 711341
                                                  30'd    8664    : data = 32'h    1D742593    ;    //    slti x11 x8 471      ====        slti a1, s0, 471
                                                  30'd    8665    : data = 32'h    41CADB33    ;    //    sra x22 x21 x28      ====        sra s6, s5, t3
                                                  30'd    8666    : data = 32'h    41FC5BB3    ;    //    sra x23 x24 x31      ====        sra s7, s8, t6
                                                  30'd    8667    : data = 32'h    01E50B33    ;    //    add x22 x10 x30      ====        add s6, a0, t5
                                                  30'd    8668    : data = 32'h    3F9BD937    ;    //    lui x18 260541      ====        lui s2, 260541
                                                  30'd    8669    : data = 32'h    00CD34B3    ;    //    sltu x9 x26 x12      ====        sltu s1, s10, a2
                                                  30'd    8670    : data = 32'h    FDB5EF93    ;    //    ori x31 x11 -37      ====        ori t6, a1, -37
                                                  30'd    8671    : data = 32'h    01B2BE33    ;    //    sltu x28 x5 x27      ====        sltu t3, t0, s11
                                                  30'd    8672    : data = 32'h    0197BC33    ;    //    sltu x24 x15 x25      ====        sltu s8, a5, s9
                                                  30'd    8673    : data = 32'h    00F592B3    ;    //    sll x5 x11 x15      ====        sll t0, a1, a5
                                                  30'd    8674    : data = 32'h    BDC6FF93    ;    //    andi x31 x13 -1060      ====        andi t6, a3, -1060
                                                  30'd    8675    : data = 32'h    72D8AD93    ;    //    slti x27 x17 1837      ====        slti s11, a7, 1837
                                                  30'd    8676    : data = 32'h    EDFA2E13    ;    //    slti x28 x20 -289      ====        slti t3, s4, -289
                                                  30'd    8677    : data = 32'h    B40E7793    ;    //    andi x15 x28 -1216      ====        andi a5, t3, -1216
                                                  30'd    8678    : data = 32'h    2329F097    ;    //    auipc x1 144031      ====        auipc ra, 144031
                                                  30'd    8679    : data = 32'h    019D2133    ;    //    slt x2 x26 x25      ====        slt sp, s10, s9
                                                  30'd    8680    : data = 32'h    014E69B3    ;    //    or x19 x28 x20      ====        or s3, t3, s4
                                                  30'd    8681    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8682    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8683    : data = 32'h    00EA16B3    ;    //    sll x13 x20 x14      ====        sll a3, s4, a4
                                                  30'd    8684    : data = 32'h    01B563B3    ;    //    or x7 x10 x27      ====        or t2, a0, s11
                                                  30'd    8685    : data = 32'h    00C05093    ;    //    srli x1 x0 12      ====        srli ra, zero, 12
                                                  30'd    8686    : data = 32'h    4031D093    ;    //    srai x1 x3 3      ====        srai ra, gp, 3
                                                  30'd    8687    : data = 32'h    E433A013    ;    //    slti x0 x7 -445      ====        slti zero, t2, -445
                                                  30'd    8688    : data = 32'h    01A8FC33    ;    //    and x24 x17 x26      ====        and s8, a7, s10
                                                  30'd    8689    : data = 32'h    00FF9CB3    ;    //    sll x25 x31 x15      ====        sll s9, t6, a5
                                                  30'd    8690    : data = 32'h    011260B3    ;    //    or x1 x4 x17      ====        or ra, tp, a7
                                                  30'd    8691    : data = 32'h    00A29E33    ;    //    sll x28 x5 x10      ====        sll t3, t0, a0
                                                  30'd    8692    : data = 32'h    00171393    ;    //    slli x7 x14 1      ====        slli t2, a4, 1
                                                  30'd    8693    : data = 32'h    30C4B713    ;    //    sltiu x14 x9 780      ====        sltiu a4, s1, 780
                                                  30'd    8694    : data = 32'h    41AA5A33    ;    //    sra x20 x20 x26      ====        sra s4, s4, s10
                                                  30'd    8695    : data = 32'h    31D12193    ;    //    slti x3 x2 797      ====        slti gp, sp, 797
                                                  30'd    8696    : data = 32'h    406E5E13    ;    //    srai x28 x28 6      ====        srai t3, t3, 6
                                                  30'd    8697    : data = 32'h    004EFD33    ;    //    and x26 x29 x4      ====        and s10, t4, tp
                                                  30'd    8698    : data = 32'h    19F3DFB7    ;    //    lui x31 106301      ====        lui t6, 106301
                                                  30'd    8699    : data = 32'h    34148F93    ;    //    addi x31 x9 833      ====        addi t6, s1, 833
                                                  30'd    8700    : data = 32'h    EE0A4313    ;    //    xori x6 x20 -288      ====        xori t1, s4, -288
                                                  30'd    8701    : data = 32'h    0AE5AD13    ;    //    slti x26 x11 174      ====        slti s10, a1, 174
                                                  30'd    8702    : data = 32'h    01385BB3    ;    //    srl x23 x16 x19      ====        srl s7, a6, s3
                                                  30'd    8703    : data = 32'h    7CFD8593    ;    //    addi x11 x27 1999      ====        addi a1, s11, 1999
                                                  30'd    8704    : data = 32'h    FBE78637    ;    //    lui x12 1031800      ====        lui a2, 1031800
                                                  30'd    8705    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8706    : data = 32'h    01D4F5B3    ;    //    and x11 x9 x29      ====        and a1, s1, t4
                                                  30'd    8707    : data = 32'h    38153113    ;    //    sltiu x2 x10 897      ====        sltiu sp, a0, 897
                                                  30'd    8708    : data = 32'h    3C193D13    ;    //    sltiu x26 x18 961      ====        sltiu s10, s2, 961
                                                  30'd    8709    : data = 32'h    01A61C93    ;    //    slli x25 x12 26      ====        slli s9, a2, 26
                                                  30'd    8710    : data = 32'h    41726D13    ;    //    ori x26 x4 1047      ====        ori s10, tp, 1047
                                                  30'd    8711    : data = 32'h    34FEEDB7    ;    //    lui x27 217070      ====        lui s11, 217070
                                                  30'd    8712    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8713    : data = 32'h    42D6B413    ;    //    sltiu x8 x13 1069      ====        sltiu s0, a3, 1069
                                                  30'd    8714    : data = 32'h    00E3CA33    ;    //    xor x20 x7 x14      ====        xor s4, t2, a4
                                                  30'd    8715    : data = 32'h    A2ADE013    ;    //    ori x0 x27 -1494      ====        ori zero, s11, -1494
                                                  30'd    8716    : data = 32'h    00767DB3    ;    //    and x27 x12 x7      ====        and s11, a2, t2
                                                  30'd    8717    : data = 32'h    00635813    ;    //    srli x16 x6 6      ====        srli a6, t1, 6
                                                  30'd    8718    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8719    : data = 32'h    22BB5717    ;    //    auipc x14 142261      ====        auipc a4, 142261
                                                  30'd    8720    : data = 32'h    0121DFB3    ;    //    srl x31 x3 x18      ====        srl t6, gp, s2
                                                  30'd    8721    : data = 32'h    00789033    ;    //    sll x0 x17 x7      ====        sll zero, a7, t2
                                                  30'd    8722    : data = 32'h    0133D093    ;    //    srli x1 x7 19      ====        srli ra, t2, 19
                                                  30'd    8723    : data = 32'h    05C2E837    ;    //    lui x16 23598      ====        lui a6, 23598
                                                  30'd    8724    : data = 32'h    4ED14BB7    ;    //    lui x23 322836      ====        lui s7, 322836
                                                  30'd    8725    : data = 32'h    41055313    ;    //    srai x6 x10 16      ====        srai t1, a0, 16
                                                  30'd    8726    : data = 32'h    00E75C13    ;    //    srli x24 x14 14      ====        srli s8, a4, 14
                                                  30'd    8727    : data = 32'h    40D4D133    ;    //    sra x2 x9 x13      ====        sra sp, s1, a3
                                                  30'd    8728    : data = 32'h    D9297C97    ;    //    auipc x25 889495      ====        auipc s9, 889495
                                                  30'd    8729    : data = 32'h    00B19A13    ;    //    slli x20 x3 11      ====        slli s4, gp, 11
                                                  30'd    8730    : data = 32'h    F971FB17    ;    //    auipc x22 1021727      ====        auipc s6, 1021727
                                                  30'd    8731    : data = 32'h    EE91C693    ;    //    xori x13 x3 -279      ====        xori a3, gp, -279
                                                  30'd    8732    : data = 32'h    002CD293    ;    //    srli x5 x25 2      ====        srli t0, s9, 2
                                                  30'd    8733    : data = 32'h    015AB333    ;    //    sltu x6 x21 x21      ====        sltu t1, s5, s5
                                                  30'd    8734    : data = 32'h    BF853293    ;    //    sltiu x5 x10 -1032      ====        sltiu t0, a0, -1032
                                                  30'd    8735    : data = 32'h    40E5DE13    ;    //    srai x28 x11 14      ====        srai t3, a1, 14
                                                  30'd    8736    : data = 32'h    F9860E93    ;    //    addi x29 x12 -104      ====        addi t4, a2, -104
                                                  30'd    8737    : data = 32'h    00EBDC93    ;    //    srli x25 x23 14      ====        srli s9, s7, 14
                                                  30'd    8738    : data = 32'h    41AD8DB3    ;    //    sub x27 x27 x26      ====        sub s11, s11, s10
                                                  30'd    8739    : data = 32'h    00DD62B3    ;    //    or x5 x26 x13      ====        or t0, s10, a3
                                                  30'd    8740    : data = 32'h    2AC10D93    ;    //    addi x27 x2 684      ====        addi s11, sp, 684
                                                  30'd    8741    : data = 32'h    00F72733    ;    //    slt x14 x14 x15      ====        slt a4, a4, a5
                                                  30'd    8742    : data = 32'h    00F89E33    ;    //    sll x28 x17 x15      ====        sll t3, a7, a5
                                                  30'd    8743    : data = 32'h    003706B3    ;    //    add x13 x14 x3      ====        add a3, a4, gp
                                                  30'd    8744    : data = 32'h    417DDDB3    ;    //    sra x27 x27 x23      ====        sra s11, s11, s7
                                                  30'd    8745    : data = 32'h    10A7CC97    ;    //    auipc x25 68220      ====        auipc s9, 68220
                                                  30'd    8746    : data = 32'h    F6C5F393    ;    //    andi x7 x11 -148      ====        andi t2, a1, -148
                                                  30'd    8747    : data = 32'h    014F6D33    ;    //    or x26 x30 x20      ====        or s10, t5, s4
                                                  30'd    8748    : data = 32'h    00A15FB3    ;    //    srl x31 x2 x10      ====        srl t6, sp, a0
                                                  30'd    8749    : data = 32'h    C7EA2713    ;    //    slti x14 x20 -898      ====        slti a4, s4, -898
                                                  30'd    8750    : data = 32'h    41378EB3    ;    //    sub x29 x15 x19      ====        sub t4, a5, s3
                                                  30'd    8751    : data = 32'h    41E35033    ;    //    sra x0 x6 x30      ====        sra zero, t1, t5
                                                  30'd    8752    : data = 32'h    3C5E0B93    ;    //    addi x23 x28 965      ====        addi s7, t3, 965
                                                  30'd    8753    : data = 32'h    E7BE0713    ;    //    addi x14 x28 -389      ====        addi a4, t3, -389
                                                  30'd    8754    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8755    : data = 32'h    6A3B2713    ;    //    slti x14 x22 1699      ====        slti a4, s6, 1699
                                                  30'd    8756    : data = 32'h    12158D37    ;    //    lui x26 74072      ====        lui s10, 74072
                                                  30'd    8757    : data = 32'h    13E8AC93    ;    //    slti x25 x17 318      ====        slti s9, a7, 318
                                                  30'd    8758    : data = 32'h    01A3D733    ;    //    srl x14 x7 x26      ====        srl a4, t2, s10
                                                  30'd    8759    : data = 32'h    000A1C13    ;    //    slli x24 x20 0      ====        slli s8, s4, 0
                                                  30'd    8760    : data = 32'h    017C1F93    ;    //    slli x31 x24 23      ====        slli t6, s8, 23
                                                  30'd    8761    : data = 32'h    01913CB3    ;    //    sltu x25 x2 x25      ====        sltu s9, sp, s9
                                                  30'd    8762    : data = 32'h    01B5E633    ;    //    or x12 x11 x27      ====        or a2, a1, s11
                                                  30'd    8763    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8764    : data = 32'h    006C65B3    ;    //    or x11 x24 x6      ====        or a1, s8, t1
                                                  30'd    8765    : data = 32'h    00C89D93    ;    //    slli x27 x17 12      ====        slli s11, a7, 12
                                                  30'd    8766    : data = 32'h    CD44AC93    ;    //    slti x25 x9 -812      ====        slti s9, s1, -812
                                                  30'd    8767    : data = 32'h    01C561B3    ;    //    or x3 x10 x28      ====        or gp, a0, t3
                                                  30'd    8768    : data = 32'h    01442FB3    ;    //    slt x31 x8 x20      ====        slt t6, s0, s4
                                                  30'd    8769    : data = 32'h    00DBB9B3    ;    //    sltu x19 x23 x13      ====        sltu s3, s7, a3
                                                  30'd    8770    : data = 32'h    FC426613    ;    //    ori x12 x4 -60      ====        ori a2, tp, -60
                                                  30'd    8771    : data = 32'h    A8ECA693    ;    //    slti x13 x25 -1394      ====        slti a3, s9, -1394
                                                  30'd    8772    : data = 32'h    B9EF4193    ;    //    xori x3 x30 -1122      ====        xori gp, t5, -1122
                                                  30'd    8773    : data = 32'h    409D84B3    ;    //    sub x9 x27 x9      ====        sub s1, s11, s1
                                                  30'd    8774    : data = 32'h    41EE03B3    ;    //    sub x7 x28 x30      ====        sub t2, t3, t5
                                                  30'd    8775    : data = 32'h    B30DEB13    ;    //    ori x22 x27 -1232      ====        ori s6, s11, -1232
                                                  30'd    8776    : data = 32'h    B5CAAE93    ;    //    slti x29 x21 -1188      ====        slti t4, s5, -1188
                                                  30'd    8777    : data = 32'h    00826A33    ;    //    or x20 x4 x8      ====        or s4, tp, s0
                                                  30'd    8778    : data = 32'h    01680333    ;    //    add x6 x16 x22      ====        add t1, a6, s6
                                                  30'd    8779    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8780    : data = 32'h    418B0333    ;    //    sub x6 x22 x24      ====        sub t1, s6, s8
                                                  30'd    8781    : data = 32'h    F31D4A93    ;    //    xori x21 x26 -207      ====        xori s5, s10, -207
                                                  30'd    8782    : data = 32'h    01152933    ;    //    slt x18 x10 x17      ====        slt s2, a0, a7
                                                  30'd    8783    : data = 32'h    41F75D33    ;    //    sra x26 x14 x31      ====        sra s10, a4, t6
                                                  30'd    8784    : data = 32'h    8F46EB93    ;    //    ori x23 x13 -1804      ====        ori s7, a3, -1804
                                                  30'd    8785    : data = 32'h    000C5E33    ;    //    srl x28 x24 x0      ====        srl t3, s8, zero
                                                  30'd    8786    : data = 32'h    00B29D93    ;    //    slli x27 x5 11      ====        slli s11, t0, 11
                                                  30'd    8787    : data = 32'h    BB603113    ;    //    sltiu x2 x0 -1098      ====        sltiu sp, zero, -1098
                                                  30'd    8788    : data = 32'h    000C2FB3    ;    //    slt x31 x24 x0      ====        slt t6, s8, zero
                                                  30'd    8789    : data = 32'h    018A7A33    ;    //    and x20 x20 x24      ====        and s4, s4, s8
                                                  30'd    8790    : data = 32'h    4008D733    ;    //    sra x14 x17 x0      ====        sra a4, a7, zero
                                                  30'd    8791    : data = 32'h    01897633    ;    //    and x12 x18 x24      ====        and a2, s2, s8
                                                  30'd    8792    : data = 32'h    00B0D793    ;    //    srli x15 x1 11      ====        srli a5, ra, 11
                                                  30'd    8793    : data = 32'h    00D53633    ;    //    sltu x12 x10 x13      ====        sltu a2, a0, a3
                                                  30'd    8794    : data = 32'h    A2886A13    ;    //    ori x20 x16 -1496      ====        ori s4, a6, -1496
                                                  30'd    8795    : data = 32'h    01BA9C93    ;    //    slli x25 x21 27      ====        slli s9, s5, 27
                                                  30'd    8796    : data = 32'h    41525893    ;    //    srai x17 x4 21      ====        srai a7, tp, 21
                                                  30'd    8797    : data = 32'h    00011833    ;    //    sll x16 x2 x0      ====        sll a6, sp, zero
                                                  30'd    8798    : data = 32'h    5E07E5B7    ;    //    lui x11 385150      ====        lui a1, 385150
                                                  30'd    8799    : data = 32'h    40A985B3    ;    //    sub x11 x19 x10      ====        sub a1, s3, a0
                                                  30'd    8800    : data = 32'h    70748793    ;    //    addi x15 x9 1799      ====        addi a5, s1, 1799
                                                  30'd    8801    : data = 32'h    0179D293    ;    //    srli x5 x19 23      ====        srli t0, s3, 23
                                                  30'd    8802    : data = 32'h    0023FC33    ;    //    and x24 x7 x2      ====        and s8, t2, sp
                                                  30'd    8803    : data = 32'h    016F0A33    ;    //    add x20 x30 x22      ====        add s4, t5, s6
                                                  30'd    8804    : data = 32'h    09416013    ;    //    ori x0 x2 148      ====        ori zero, sp, 148
                                                  30'd    8805    : data = 32'h    005F4633    ;    //    xor x12 x30 x5      ====        xor a2, t5, t0
                                                  30'd    8806    : data = 32'h    01B6F333    ;    //    and x6 x13 x27      ====        and t1, a3, s11
                                                  30'd    8807    : data = 32'h    0D628037    ;    //    lui x0 54824      ====        lui zero, 54824
                                                  30'd    8808    : data = 32'h    7E5F4D93    ;    //    xori x27 x30 2021      ====        xori s11, t5, 2021
                                                  30'd    8809    : data = 32'h    413E51B3    ;    //    sra x3 x28 x19      ====        sra gp, t3, s3
                                                  30'd    8810    : data = 32'h    4EBDB393    ;    //    sltiu x7 x27 1259      ====        sltiu t2, s11, 1259
                                                  30'd    8811    : data = 32'h    01F41FB3    ;    //    sll x31 x8 x31      ====        sll t6, s0, t6
                                                  30'd    8812    : data = 32'h    EDD37913    ;    //    andi x18 x6 -291      ====        andi s2, t1, -291
                                                  30'd    8813    : data = 32'h    01982B13    ;    //    slti x22 x16 25      ====        slti s6, a6, 25
                                                  30'd    8814    : data = 32'h    01049713    ;    //    slli x14 x9 16      ====        slli a4, s1, 16
                                                  30'd    8815    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8816    : data = 32'h    4026DE13    ;    //    srai x28 x13 2      ====        srai t3, a3, 2
                                                  30'd    8817    : data = 32'h    3ECBCA13    ;    //    xori x20 x23 1004      ====        xori s4, s7, 1004
                                                  30'd    8818    : data = 32'h    001F5C13    ;    //    srli x24 x30 1      ====        srli s8, t5, 1
                                                  30'd    8819    : data = 32'h    A9BB0593    ;    //    addi x11 x22 -1381      ====        addi a1, s6, -1381
                                                  30'd    8820    : data = 32'h    000B9BB3    ;    //    sll x23 x23 x0      ====        sll s7, s7, zero
                                                  30'd    8821    : data = 32'h    222D2D13    ;    //    slti x26 x26 546      ====        slti s10, s10, 546
                                                  30'd    8822    : data = 32'h    41890E33    ;    //    sub x28 x18 x24      ====        sub t3, s2, s8
                                                  30'd    8823    : data = 32'h    AB760F93    ;    //    addi x31 x12 -1353      ====        addi t6, a2, -1353
                                                  30'd    8824    : data = 32'h    90F24313    ;    //    xori x6 x4 -1777      ====        xori t1, tp, -1777
                                                  30'd    8825    : data = 32'h    00880D33    ;    //    add x26 x16 x8      ====        add s10, a6, s0
                                                  30'd    8826    : data = 32'h    0130DD93    ;    //    srli x27 x1 19      ====        srli s11, ra, 19
                                                  30'd    8827    : data = 32'h    F36EBCB7    ;    //    lui x25 997099      ====        lui s9, 997099
                                                  30'd    8828    : data = 32'h    413F5033    ;    //    sra x0 x30 x19      ====        sra zero, t5, s3
                                                  30'd    8829    : data = 32'h    01102733    ;    //    slt x14 x0 x17      ====        slt a4, zero, a7
                                                  30'd    8830    : data = 32'h    01C87C33    ;    //    and x24 x16 x28      ====        and s8, a6, t3
                                                  30'd    8831    : data = 32'h    01AC9CB3    ;    //    sll x25 x25 x26      ====        sll s9, s9, s10
                                                  30'd    8832    : data = 32'h    013E5113    ;    //    srli x2 x28 19      ====        srli sp, t3, 19
                                                  30'd    8833    : data = 32'h    01793BB3    ;    //    sltu x23 x18 x23      ====        sltu s7, s2, s7
                                                  30'd    8834    : data = 32'h    74CA3B93    ;    //    sltiu x23 x20 1868      ====        sltiu s7, s4, 1868
                                                  30'd    8835    : data = 32'h    D9E7E493    ;    //    ori x9 x15 -610      ====        ori s1, a5, -610
                                                  30'd    8836    : data = 32'h    002C7833    ;    //    and x16 x24 x2      ====        and a6, s8, sp
                                                  30'd    8837    : data = 32'h    79A7EC13    ;    //    ori x24 x15 1946      ====        ori s8, a5, 1946
                                                  30'd    8838    : data = 32'h    322FBE13    ;    //    sltiu x28 x31 802      ====        sltiu t3, t6, 802
                                                  30'd    8839    : data = 32'h    00611013    ;    //    slli x0 x2 6      ====        slli zero, sp, 6
                                                  30'd    8840    : data = 32'h    006AB633    ;    //    sltu x12 x21 x6      ====        sltu a2, s5, t1
                                                  30'd    8841    : data = 32'h    00F85733    ;    //    srl x14 x16 x15      ====        srl a4, a6, a5
                                                  30'd    8842    : data = 32'h    4D9A2C93    ;    //    slti x25 x20 1241      ====        slti s9, s4, 1241
                                                  30'd    8843    : data = 32'h    14B0F897    ;    //    auipc x17 84751      ====        auipc a7, 84751
                                                  30'd    8844    : data = 32'h    1E0A0713    ;    //    addi x14 x20 480      ====        addi a4, s4, 480
                                                  30'd    8845    : data = 32'h    005FCC33    ;    //    xor x24 x31 x5      ====        xor s8, t6, t0
                                                  30'd    8846    : data = 32'h    00D1DB93    ;    //    srli x23 x3 13      ====        srli s7, gp, 13
                                                  30'd    8847    : data = 32'h    00289A93    ;    //    slli x21 x17 2      ====        slli s5, a7, 2
                                                  30'd    8848    : data = 32'h    01C3CE33    ;    //    xor x28 x7 x28      ====        xor t3, t2, t3
                                                  30'd    8849    : data = 32'h    0194DC33    ;    //    srl x24 x9 x25      ====        srl s8, s1, s9
                                                  30'd    8850    : data = 32'h    410580B3    ;    //    sub x1 x11 x16      ====        sub ra, a1, a6
                                                  30'd    8851    : data = 32'h    4109D113    ;    //    srai x2 x19 16      ====        srai sp, s3, 16
                                                  30'd    8852    : data = 32'h    01BC5113    ;    //    srli x2 x24 27      ====        srli sp, s8, 27
                                                  30'd    8853    : data = 32'h    01B54833    ;    //    xor x16 x10 x27      ====        xor a6, a0, s11
                                                  30'd    8854    : data = 32'h    014B68B3    ;    //    or x17 x22 x20      ====        or a7, s6, s4
                                                  30'd    8855    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8856    : data = 32'h    00B29813    ;    //    slli x16 x5 11      ====        slli a6, t0, 11
                                                  30'd    8857    : data = 32'h    0032DD13    ;    //    srli x26 x5 3      ====        srli s10, t0, 3
                                                  30'd    8858    : data = 32'h    41865B93    ;    //    srai x23 x12 24      ====        srai s7, a2, 24
                                                  30'd    8859    : data = 32'h    008AAC33    ;    //    slt x24 x21 x8      ====        slt s8, s5, s0
                                                  30'd    8860    : data = 32'h    01577833    ;    //    and x16 x14 x21      ====        and a6, a4, s5
                                                  30'd    8861    : data = 32'h    E57D0493    ;    //    addi x9 x26 -425      ====        addi s1, s10, -425
                                                  30'd    8862    : data = 32'h    01C73BB3    ;    //    sltu x23 x14 x28      ====        sltu s7, a4, t3
                                                  30'd    8863    : data = 32'h    013455B3    ;    //    srl x11 x8 x19      ====        srl a1, s0, s3
                                                  30'd    8864    : data = 32'h    019D9A13    ;    //    slli x20 x27 25      ====        slli s4, s11, 25
                                                  30'd    8865    : data = 32'h    016B9D93    ;    //    slli x27 x23 22      ====        slli s11, s7, 22
                                                  30'd    8866    : data = 32'h    01D51333    ;    //    sll x6 x10 x29      ====        sll t1, a0, t4
                                                  30'd    8867    : data = 32'h    041B0793    ;    //    addi x15 x22 65      ====        addi a5, s6, 65
                                                  30'd    8868    : data = 32'h    017905B3    ;    //    add x11 x18 x23      ====        add a1, s2, s7
                                                  30'd    8869    : data = 32'h    0169D333    ;    //    srl x6 x19 x22      ====        srl t1, s3, s6
                                                  30'd    8870    : data = 32'h    41B7DFB3    ;    //    sra x31 x15 x27      ====        sra t6, a5, s11
                                                  30'd    8871    : data = 32'h    40FB8A33    ;    //    sub x20 x23 x15      ====        sub s4, s7, a5
                                                  30'd    8872    : data = 32'h    A763AD13    ;    //    slti x26 x7 -1418      ====        slti s10, t2, -1418
                                                  30'd    8873    : data = 32'h    00211C33    ;    //    sll x24 x2 x2      ====        sll s8, sp, sp
                                                  30'd    8874    : data = 32'h    0116B8B3    ;    //    sltu x17 x13 x17      ====        sltu a7, a3, a7
                                                  30'd    8875    : data = 32'h    01789393    ;    //    slli x7 x17 23      ====        slli t2, a7, 23
                                                  30'd    8876    : data = 32'h    004664B3    ;    //    or x9 x12 x4      ====        or s1, a2, tp
                                                  30'd    8877    : data = 32'h    00717833    ;    //    and x16 x2 x7      ====        and a6, sp, t2
                                                  30'd    8878    : data = 32'h    E9EEC613    ;    //    xori x12 x29 -354      ====        xori a2, t4, -354
                                                  30'd    8879    : data = 32'h    417052B3    ;    //    sra x5 x0 x23      ====        sra t0, zero, s7
                                                  30'd    8880    : data = 32'h    01099633    ;    //    sll x12 x19 x16      ====        sll a2, s3, a6
                                                  30'd    8881    : data = 32'h    D0F6C813    ;    //    xori x16 x13 -753      ====        xori a6, a3, -753
                                                  30'd    8882    : data = 32'h    C7F24B93    ;    //    xori x23 x4 -897      ====        xori s7, tp, -897
                                                  30'd    8883    : data = 32'h    00D64833    ;    //    xor x16 x12 x13      ====        xor a6, a2, a3
                                                  30'd    8884    : data = 32'h    002967B3    ;    //    or x15 x18 x2      ====        or a5, s2, sp
                                                  30'd    8885    : data = 32'h    001697B3    ;    //    sll x15 x13 x1      ====        sll a5, a3, ra
                                                  30'd    8886    : data = 32'h    008A6D33    ;    //    or x26 x20 x8      ====        or s10, s4, s0
                                                  30'd    8887    : data = 32'h    82B40B37    ;    //    lui x22 535360      ====        lui s6, 535360
                                                  30'd    8888    : data = 32'h    40725D13    ;    //    srai x26 x4 7      ====        srai s10, tp, 7
                                                  30'd    8889    : data = 32'h    09ACB993    ;    //    sltiu x19 x25 154      ====        sltiu s3, s9, 154
                                                  30'd    8890    : data = 32'h    00DBEB33    ;    //    or x22 x23 x13      ====        or s6, s7, a3
                                                  30'd    8891    : data = 32'h    077EBC13    ;    //    sltiu x24 x29 119      ====        sltiu s8, t4, 119
                                                  30'd    8892    : data = 32'h    0F61BA93    ;    //    sltiu x21 x3 246      ====        sltiu s5, gp, 246
                                                  30'd    8893    : data = 32'h    01D2DC33    ;    //    srl x24 x5 x29      ====        srl s8, t0, t4
                                                  30'd    8894    : data = 32'h    006445B3    ;    //    xor x11 x8 x6      ====        xor a1, s0, t1
                                                  30'd    8895    : data = 32'h    001DC2B3    ;    //    xor x5 x27 x1      ====        xor t0, s11, ra
                                                  30'd    8896    : data = 32'h    41B4D013    ;    //    srai x0 x9 27      ====        srai zero, s1, 27
                                                  30'd    8897    : data = 32'h    3DD52437    ;    //    lui x8 253266      ====        lui s0, 253266
                                                  30'd    8898    : data = 32'h    01690433    ;    //    add x8 x18 x22      ====        add s0, s2, s6
                                                  30'd    8899    : data = 32'h    934FCA93    ;    //    xori x21 x31 -1740      ====        xori s5, t6, -1740
                                                  30'd    8900    : data = 32'h    9CB7B013    ;    //    sltiu x0 x15 -1589      ====        sltiu zero, a5, -1589
                                                  30'd    8901    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8902    : data = 32'h    401A5093    ;    //    srai x1 x20 1      ====        srai ra, s4, 1
                                                  30'd    8903    : data = 32'h    55E20D13    ;    //    addi x26 x4 1374      ====        addi s10, tp, 1374
                                                  30'd    8904    : data = 32'h    0AEA0713    ;    //    addi x14 x20 174      ====        addi a4, s4, 174
                                                  30'd    8905    : data = 32'h    004DBB33    ;    //    sltu x22 x27 x4      ====        sltu s6, s11, tp
                                                  30'd    8906    : data = 32'h    00CB9D13    ;    //    slli x26 x23 12      ====        slli s10, s7, 12
                                                  30'd    8907    : data = 32'h    73A36693    ;    //    ori x13 x6 1850      ====        ori a3, t1, 1850
                                                  30'd    8908    : data = 32'h    401D0C33    ;    //    sub x24 x26 x1      ====        sub s8, s10, ra
                                                  30'd    8909    : data = 32'h    418E5193    ;    //    srai x3 x28 24      ====        srai gp, t3, 24
                                                  30'd    8910    : data = 32'h    009C58B3    ;    //    srl x17 x24 x9      ====        srl a7, s8, s1
                                                  30'd    8911    : data = 32'h    A8AC8C37    ;    //    lui x24 690888      ====        lui s8, 690888
                                                  30'd    8912    : data = 32'h    00511193    ;    //    slli x3 x2 5      ====        slli gp, sp, 5
                                                  30'd    8913    : data = 32'h    30CEAC13    ;    //    slti x24 x29 780      ====        slti s8, t4, 780
                                                  30'd    8914    : data = 32'h    01133033    ;    //    sltu x0 x6 x17      ====        sltu zero, t1, a7
                                                  30'd    8915    : data = 32'h    0187C1B3    ;    //    xor x3 x15 x24      ====        xor gp, a5, s8
                                                  30'd    8916    : data = 32'h    76AC2017    ;    //    auipc x0 486082      ====        auipc zero, 486082
                                                  30'd    8917    : data = 32'h    00E02933    ;    //    slt x18 x0 x14      ====        slt s2, zero, a4
                                                  30'd    8918    : data = 32'h    22D7F113    ;    //    andi x2 x15 557      ====        andi sp, a5, 557
                                                  30'd    8919    : data = 32'h    74DA7293    ;    //    andi x5 x20 1869      ====        andi t0, s4, 1869
                                                  30'd    8920    : data = 32'h    B8EEBA13    ;    //    sltiu x20 x29 -1138      ====        sltiu s4, t4, -1138
                                                  30'd    8921    : data = 32'h    00955793    ;    //    srli x15 x10 9      ====        srli a5, a0, 9
                                                  30'd    8922    : data = 32'h    01F7FC33    ;    //    and x24 x15 x31      ====        and s8, a5, t6
                                                  30'd    8923    : data = 32'h    13F68713    ;    //    addi x14 x13 319      ====        addi a4, a3, 319
                                                  30'd    8924    : data = 32'h    4188D633    ;    //    sra x12 x17 x24      ====        sra a2, a7, s8
                                                  30'd    8925    : data = 32'h    0D8025B7    ;    //    lui x11 55298      ====        lui a1, 55298
                                                  30'd    8926    : data = 32'h    59493813    ;    //    sltiu x16 x18 1428      ====        sltiu a6, s2, 1428
                                                  30'd    8927    : data = 32'h    A40BCDB7    ;    //    lui x27 671932      ====        lui s11, 671932
                                                  30'd    8928    : data = 32'h    01F91293    ;    //    slli x5 x18 31      ====        slli t0, s2, 31
                                                  30'd    8929    : data = 32'h    90E87093    ;    //    andi x1 x16 -1778      ====        andi ra, a6, -1778
                                                  30'd    8930    : data = 32'h    01C4FCB3    ;    //    and x25 x9 x28      ====        and s9, s1, t3
                                                  30'd    8931    : data = 32'h    0139F933    ;    //    and x18 x19 x19      ====        and s2, s3, s3
                                                  30'd    8932    : data = 32'h    F1286F93    ;    //    ori x31 x16 -238      ====        ori t6, a6, -238
                                                  30'd    8933    : data = 32'h    D2D9CA13    ;    //    xori x20 x19 -723      ====        xori s4, s3, -723
                                                  30'd    8934    : data = 32'h    B1A46137    ;    //    lui x2 727622      ====        lui sp, 727622
                                                  30'd    8935    : data = 32'h    A3A27693    ;    //    andi x13 x4 -1478      ====        andi a3, tp, -1478
                                                  30'd    8936    : data = 32'h    003FBC33    ;    //    sltu x24 x31 x3      ====        sltu s8, t6, gp
                                                  30'd    8937    : data = 32'h    00D3CD33    ;    //    xor x26 x7 x13      ====        xor s10, t2, a3
                                                  30'd    8938    : data = 32'h    41168D33    ;    //    sub x26 x13 x17      ====        sub s10, a3, a7
                                                  30'd    8939    : data = 32'h    017CF033    ;    //    and x0 x25 x23      ====        and zero, s9, s7
                                                  30'd    8940    : data = 32'h    012165B3    ;    //    or x11 x2 x18      ====        or a1, sp, s2
                                                  30'd    8941    : data = 32'h    40A3DC33    ;    //    sra x24 x7 x10      ====        sra s8, t2, a0
                                                  30'd    8942    : data = 32'h    01D3E2B3    ;    //    or x5 x7 x29      ====        or t0, t2, t4
                                                  30'd    8943    : data = 32'h    9B4ABA13    ;    //    sltiu x20 x21 -1612      ====        sltiu s4, s5, -1612
                                                  30'd    8944    : data = 32'h    7B54E093    ;    //    ori x1 x9 1973      ====        ori ra, s1, 1973
                                                  30'd    8945    : data = 32'h    014334B3    ;    //    sltu x9 x6 x20      ====        sltu s1, t1, s4
                                                  30'd    8946    : data = 32'h    EF0F3593    ;    //    sltiu x11 x30 -272      ====        sltiu a1, t5, -272
                                                  30'd    8947    : data = 32'h    40AD0AB3    ;    //    sub x21 x26 x10      ====        sub s5, s10, a0
                                                  30'd    8948    : data = 32'h    01C3B033    ;    //    sltu x0 x7 x28      ====        sltu zero, t2, t3
                                                  30'd    8949    : data = 32'h    002DF433    ;    //    and x8 x27 x2      ====        and s0, s11, sp
                                                  30'd    8950    : data = 32'h    40B309B3    ;    //    sub x19 x6 x11      ====        sub s3, t1, a1
                                                  30'd    8951    : data = 32'h    F007BE13    ;    //    sltiu x28 x15 -256      ====        sltiu t3, a5, -256
                                                  30'd    8952    : data = 32'h    0098CB33    ;    //    xor x22 x17 x9      ====        xor s6, a7, s1
                                                  30'd    8953    : data = 32'h    00241E93    ;    //    slli x29 x8 2      ====        slli t4, s0, 2
                                                  30'd    8954    : data = 32'h    00FCDD93    ;    //    srli x27 x25 15      ====        srli s11, s9, 15
                                                  30'd    8955    : data = 32'h    40B75193    ;    //    srai x3 x14 11      ====        srai gp, a4, 11
                                                  30'd    8956    : data = 32'h    41BF5D93    ;    //    srai x27 x30 27      ====        srai s11, t5, 27
                                                  30'd    8957    : data = 32'h    E06AC637    ;    //    lui x12 919212      ====        lui a2, 919212
                                                  30'd    8958    : data = 32'h    01A87433    ;    //    and x8 x16 x26      ====        and s0, a6, s10
                                                  30'd    8959    : data = 32'h    1950E437    ;    //    lui x8 103694      ====        lui s0, 103694
                                                  30'd    8960    : data = 32'h    411552B3    ;    //    sra x5 x10 x17      ====        sra t0, a0, a7
                                                  30'd    8961    : data = 32'h    4CD8E093    ;    //    ori x1 x17 1229      ====        ori ra, a7, 1229
                                                  30'd    8962    : data = 32'h    8B49A013    ;    //    slti x0 x19 -1868      ====        slti zero, s3, -1868
                                                  30'd    8963    : data = 32'h    0022CFB3    ;    //    xor x31 x5 x2      ====        xor t6, t0, sp
                                                  30'd    8964    : data = 32'h    0044B1B3    ;    //    sltu x3 x9 x4      ====        sltu gp, s1, tp
                                                  30'd    8965    : data = 32'h    40425EB3    ;    //    sra x29 x4 x4      ====        sra t4, tp, tp
                                                  30'd    8966    : data = 32'h    6ED00C97    ;    //    auipc x25 453888      ====        auipc s9, 453888
                                                  30'd    8967    : data = 32'h    408E5033    ;    //    sra x0 x28 x8      ====        sra zero, t3, s0
                                                  30'd    8968    : data = 32'h    C4A00A13    ;    //    addi x20 x0 -950      ====        addi s4, zero, -950
                                                  30'd    8969    : data = 32'h    3CCF6D13    ;    //    ori x26 x30 972      ====        ori s10, t5, 972
                                                  30'd    8970    : data = 32'h    00FAA733    ;    //    slt x14 x21 x15      ====        slt a4, s5, a5
                                                  30'd    8971    : data = 32'h    04127913    ;    //    andi x18 x4 65      ====        andi s2, tp, 65
                                                  30'd    8972    : data = 32'h    00A68A33    ;    //    add x20 x13 x10      ====        add s4, a3, a0
                                                  30'd    8973    : data = 32'h    01CA5A33    ;    //    srl x20 x20 x28      ====        srl s4, s4, t3
                                                  30'd    8974    : data = 32'h    BB910637    ;    //    lui x12 768272      ====        lui a2, 768272
                                                  30'd    8975    : data = 32'h    30D69597    ;    //    auipc x11 200041      ====        auipc a1, 200041
                                                  30'd    8976    : data = 32'h    01C83FB3    ;    //    sltu x31 x16 x28      ====        sltu t6, a6, t3
                                                  30'd    8977    : data = 32'h    22B26D13    ;    //    ori x26 x4 555      ====        ori s10, tp, 555
                                                  30'd    8978    : data = 32'h    91D62693    ;    //    slti x13 x12 -1763      ====        slti a3, a2, -1763
                                                  30'd    8979    : data = 32'h    4019D333    ;    //    sra x6 x19 x1      ====        sra t1, s3, ra
                                                  30'd    8980    : data = 32'h    0166B133    ;    //    sltu x2 x13 x22      ====        sltu sp, a3, s6
                                                  30'd    8981    : data = 32'h    BDC98093    ;    //    addi x1 x19 -1060      ====        addi ra, s3, -1060
                                                  30'd    8982    : data = 32'h    00447FB3    ;    //    and x31 x8 x4      ====        and t6, s0, tp
                                                  30'd    8983    : data = 32'h    41EA5933    ;    //    sra x18 x20 x30      ====        sra s2, s4, t5
                                                  30'd    8984    : data = 32'h    00D29B33    ;    //    sll x22 x5 x13      ====        sll s6, t0, a3
                                                  30'd    8985    : data = 32'h    007E88B3    ;    //    add x17 x29 x7      ====        add a7, t4, t2
                                                  30'd    8986    : data = 32'h    41965733    ;    //    sra x14 x12 x25      ====        sra a4, a2, s9
                                                  30'd    8987    : data = 32'h    0100D593    ;    //    srli x11 x1 16      ====        srli a1, ra, 16
                                                  30'd    8988    : data = 32'h    C9EC2697    ;    //    auipc x13 827074      ====        auipc a3, 827074
                                                  30'd    8989    : data = 32'h    01081D33    ;    //    sll x26 x16 x16      ====        sll s10, a6, a6
                                                  30'd    8990    : data = 32'h    018FEAB3    ;    //    or x21 x31 x24      ====        or s5, t6, s8
                                                  30'd    8991    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8992    : data = 32'h    00E61613    ;    //    slli x12 x12 14      ====        slli a2, a2, 14
                                                  30'd    8993    : data = 32'h    015E0CB3    ;    //    add x25 x28 x21      ====        add s9, t3, s5
                                                  30'd    8994    : data = 32'h    DBE7EB13    ;    //    ori x22 x15 -578      ====        ori s6, a5, -578
                                                  30'd    8995    : data = 32'h    005E4B33    ;    //    xor x22 x28 x5      ====        xor s6, t3, t0
                                                  30'd    8996    : data = 32'h    1702C113    ;    //    xori x2 x5 368      ====        xori sp, t0, 368
                                                  30'd    8997    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    8998    : data = 32'h    40D20BB3    ;    //    sub x23 x4 x13      ====        sub s7, tp, a3
                                                  30'd    8999    : data = 32'h    DFE9BB37    ;    //    lui x22 917147      ====        lui s6, 917147
                                                  30'd    9000    : data = 32'h    78CBC493    ;    //    xori x9 x23 1932      ====        xori s1, s7, 1932
                                                  30'd    9001    : data = 32'h    A64232B7    ;    //    lui x5 680995      ====        lui t0, 680995
                                                  30'd    9002    : data = 32'h    018A6633    ;    //    or x12 x20 x24      ====        or a2, s4, s8
                                                  30'd    9003    : data = 32'h    BF50F013    ;    //    andi x0 x1 -1035      ====        andi zero, ra, -1035
                                                  30'd    9004    : data = 32'h    0095EAB3    ;    //    or x21 x11 x9      ====        or s5, a1, s1
                                                  30'd    9005    : data = 32'h    40858133    ;    //    sub x2 x11 x8      ====        sub sp, a1, s0
                                                  30'd    9006    : data = 32'h    0118B433    ;    //    sltu x8 x17 x17      ====        sltu s0, a7, a7
                                                  30'd    9007    : data = 32'h    C10EC613    ;    //    xori x12 x29 -1008      ====        xori a2, t4, -1008
                                                  30'd    9008    : data = 32'h    41365013    ;    //    srai x0 x12 19      ====        srai zero, a2, 19
                                                  30'd    9009    : data = 32'h    018BD9B3    ;    //    srl x19 x23 x24      ====        srl s3, s7, s8
                                                  30'd    9010    : data = 32'h    012EE333    ;    //    or x6 x29 x18      ====        or t1, t4, s2
                                                  30'd    9011    : data = 32'h    01EEDF93    ;    //    srli x31 x29 30      ====        srli t6, t4, 30
                                                  30'd    9012    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9013    : data = 32'h    003A02B3    ;    //    add x5 x20 x3      ====        add t0, s4, gp
                                                  30'd    9014    : data = 32'h    898C3D13    ;    //    sltiu x26 x24 -1896      ====        sltiu s10, s8, -1896
                                                  30'd    9015    : data = 32'h    40E7D613    ;    //    srai x12 x15 14      ====        srai a2, a5, 14
                                                  30'd    9016    : data = 32'h    014D13B3    ;    //    sll x7 x26 x20      ====        sll t2, s10, s4
                                                  30'd    9017    : data = 32'h    018910B3    ;    //    sll x1 x18 x24      ====        sll ra, s2, s8
                                                  30'd    9018    : data = 32'h    00321313    ;    //    slli x6 x4 3      ====        slli t1, tp, 3
                                                  30'd    9019    : data = 32'h    EC0BFC13    ;    //    andi x24 x23 -320      ====        andi s8, s7, -320
                                                  30'd    9020    : data = 32'h    400E5C33    ;    //    sra x24 x28 x0      ====        sra s8, t3, zero
                                                  30'd    9021    : data = 32'h    01EC08B3    ;    //    add x17 x24 x30      ====        add a7, s8, t5
                                                  30'd    9022    : data = 32'h    003A5E33    ;    //    srl x28 x20 x3      ====        srl t3, s4, gp
                                                  30'd    9023    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9024    : data = 32'h    AACF0913    ;    //    addi x18 x30 -1364      ====        addi s2, t5, -1364
                                                  30'd    9025    : data = 32'h    405D5093    ;    //    srai x1 x26 5      ====        srai ra, s10, 5
                                                  30'd    9026    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9027    : data = 32'h    00FEB4B3    ;    //    sltu x9 x29 x15      ====        sltu s1, t4, a5
                                                  30'd    9028    : data = 32'h    00CBAD33    ;    //    slt x26 x23 x12      ====        slt s10, s7, a2
                                                  30'd    9029    : data = 32'h    DB569317    ;    //    auipc x6 898409      ====        auipc t1, 898409
                                                  30'd    9030    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9031    : data = 32'h    012B2E33    ;    //    slt x28 x22 x18      ====        slt t3, s6, s2
                                                  30'd    9032    : data = 32'h    000522B3    ;    //    slt x5 x10 x0      ====        slt t0, a0, zero
                                                  30'd    9033    : data = 32'h    41D003B3    ;    //    sub x7 x0 x29      ====        sub t2, zero, t4
                                                  30'd    9034    : data = 32'h    E1285997    ;    //    auipc x19 922245      ====        auipc s3, 922245
                                                  30'd    9035    : data = 32'h    C792C613    ;    //    xori x12 x5 -903      ====        xori a2, t0, -903
                                                  30'd    9036    : data = 32'h    1BBD7093    ;    //    andi x1 x26 443      ====        andi ra, s10, 443
                                                  30'd    9037    : data = 32'h    41285A13    ;    //    srai x20 x16 18      ====        srai s4, a6, 18
                                                  30'd    9038    : data = 32'h    41585B93    ;    //    srai x23 x16 21      ====        srai s7, a6, 21
                                                  30'd    9039    : data = 32'h    01A29633    ;    //    sll x12 x5 x26      ====        sll a2, t0, s10
                                                  30'd    9040    : data = 32'h    001BC133    ;    //    xor x2 x23 x1      ====        xor sp, s7, ra
                                                  30'd    9041    : data = 32'h    516EAB93    ;    //    slti x23 x29 1302      ====        slti s7, t4, 1302
                                                  30'd    9042    : data = 32'h    0085D593    ;    //    srli x11 x11 8      ====        srli a1, a1, 8
                                                  30'd    9043    : data = 32'h    00B6A433    ;    //    slt x8 x13 x11      ====        slt s0, a3, a1
                                                  30'd    9044    : data = 32'h    0134B4B3    ;    //    sltu x9 x9 x19      ====        sltu s1, s1, s3
                                                  30'd    9045    : data = 32'h    D56FEB13    ;    //    ori x22 x31 -682      ====        ori s6, t6, -682
                                                  30'd    9046    : data = 32'h    00E86733    ;    //    or x14 x16 x14      ====        or a4, a6, a4
                                                  30'd    9047    : data = 32'h    01AC3D33    ;    //    sltu x26 x24 x26      ====        sltu s10, s8, s10
                                                  30'd    9048    : data = 32'h    002CBB33    ;    //    sltu x22 x25 x2      ====        sltu s6, s9, sp
                                                  30'd    9049    : data = 32'h    194DDB97    ;    //    auipc x23 103645      ====        auipc s7, 103645
                                                  30'd    9050    : data = 32'h    57633B93    ;    //    sltiu x23 x6 1398      ====        sltiu s7, t1, 1398
                                                  30'd    9051    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9052    : data = 32'h    003A65B3    ;    //    or x11 x20 x3      ====        or a1, s4, gp
                                                  30'd    9053    : data = 32'h    40605B93    ;    //    srai x23 x0 6      ====        srai s7, zero, 6
                                                  30'd    9054    : data = 32'h    9270BD13    ;    //    sltiu x26 x1 -1753      ====        sltiu s10, ra, -1753
                                                  30'd    9055    : data = 32'h    57C18E13    ;    //    addi x28 x3 1404      ====        addi t3, gp, 1404
                                                  30'd    9056    : data = 32'h    4034DAB3    ;    //    sra x21 x9 x3      ====        sra s5, s1, gp
                                                  30'd    9057    : data = 32'h    401185B3    ;    //    sub x11 x3 x1      ====        sub a1, gp, ra
                                                  30'd    9058    : data = 32'h    009C0D33    ;    //    add x26 x24 x9      ====        add s10, s8, s1
                                                  30'd    9059    : data = 32'h    017CC4B3    ;    //    xor x9 x25 x23      ====        xor s1, s9, s7
                                                  30'd    9060    : data = 32'h    1E016413    ;    //    ori x8 x2 480      ====        ori s0, sp, 480
                                                  30'd    9061    : data = 32'h    21317693    ;    //    andi x13 x2 531      ====        andi a3, sp, 531
                                                  30'd    9062    : data = 32'h    01ED5F93    ;    //    srli x31 x26 30      ====        srli t6, s10, 30
                                                  30'd    9063    : data = 32'h    AB0AC693    ;    //    xori x13 x21 -1360      ====        xori a3, s5, -1360
                                                  30'd    9064    : data = 32'h    001D5D13    ;    //    srli x26 x26 1      ====        srli s10, s10, 1
                                                  30'd    9065    : data = 32'h    00599033    ;    //    sll x0 x19 x5      ====        sll zero, s3, t0
                                                  30'd    9066    : data = 32'h    E8AFB413    ;    //    sltiu x8 x31 -374      ====        sltiu s0, t6, -374
                                                  30'd    9067    : data = 32'h    E3C04D93    ;    //    xori x27 x0 -452      ====        xori s11, zero, -452
                                                  30'd    9068    : data = 32'h    944E4C13    ;    //    xori x24 x28 -1724      ====        xori s8, t3, -1724
                                                  30'd    9069    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9070    : data = 32'h    B0CD69B7    ;    //    lui x19 724182      ====        lui s3, 724182
                                                  30'd    9071    : data = 32'h    4090D633    ;    //    sra x12 x1 x9      ====        sra a2, ra, s1
                                                  30'd    9072    : data = 32'h    003DD333    ;    //    srl x6 x27 x3      ====        srl t1, s11, gp
                                                  30'd    9073    : data = 32'h    271C0993    ;    //    addi x19 x24 625      ====        addi s3, s8, 625
                                                  30'd    9074    : data = 32'h    7C7BCE93    ;    //    xori x29 x23 1991      ====        xori t4, s7, 1991
                                                  30'd    9075    : data = 32'h    A7B1FD93    ;    //    andi x27 x3 -1413      ====        andi s11, gp, -1413
                                                  30'd    9076    : data = 32'h    00E7E2B3    ;    //    or x5 x15 x14      ====        or t0, a5, a4
                                                  30'd    9077    : data = 32'h    1F68E193    ;    //    ori x3 x17 502      ====        ori gp, a7, 502
                                                  30'd    9078    : data = 32'h    01BFBC33    ;    //    sltu x24 x31 x27      ====        sltu s8, t6, s11
                                                  30'd    9079    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9080    : data = 32'h    40B5D413    ;    //    srai x8 x11 11      ====        srai s0, a1, 11
                                                  30'd    9081    : data = 32'h    E23F0B13    ;    //    addi x22 x30 -477      ====        addi s6, t5, -477
                                                  30'd    9082    : data = 32'h    29E80D13    ;    //    addi x26 x16 670      ====        addi s10, a6, 670
                                                  30'd    9083    : data = 32'h    09BA2F93    ;    //    slti x31 x20 155      ====        slti t6, s4, 155
                                                  30'd    9084    : data = 32'h    409050B3    ;    //    sra x1 x0 x9      ====        sra ra, zero, s1
                                                  30'd    9085    : data = 32'h    8020E993    ;    //    ori x19 x1 -2046      ====        ori s3, ra, -2046
                                                  30'd    9086    : data = 32'h    003E4933    ;    //    xor x18 x28 x3      ====        xor s2, t3, gp
                                                  30'd    9087    : data = 32'h    00F1EE33    ;    //    or x28 x3 x15      ====        or t3, gp, a5
                                                  30'd    9088    : data = 32'h    019550B3    ;    //    srl x1 x10 x25      ====        srl ra, a0, s9
                                                  30'd    9089    : data = 32'h    015D3B33    ;    //    sltu x22 x26 x21      ====        sltu s6, s10, s5
                                                  30'd    9090    : data = 32'h    8993C293    ;    //    xori x5 x7 -1895      ====        xori t0, t2, -1895
                                                  30'd    9091    : data = 32'h    189AB713    ;    //    sltiu x14 x21 393      ====        sltiu a4, s5, 393
                                                  30'd    9092    : data = 32'h    4044DCB3    ;    //    sra x25 x9 x4      ====        sra s9, s1, tp
                                                  30'd    9093    : data = 32'h    1C655397    ;    //    auipc x7 116309      ====        auipc t2, 116309
                                                  30'd    9094    : data = 32'h    4070DBB3    ;    //    sra x23 x1 x7      ====        sra s7, ra, t2
                                                  30'd    9095    : data = 32'h    A401C013    ;    //    xori x0 x3 -1472      ====        xori zero, gp, -1472
                                                  30'd    9096    : data = 32'h    9136A013    ;    //    slti x0 x13 -1773      ====        slti zero, a3, -1773
                                                  30'd    9097    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9098    : data = 32'h    4A68EA13    ;    //    ori x20 x17 1190      ====        ori s4, a7, 1190
                                                  30'd    9099    : data = 32'h    41A6D413    ;    //    srai x8 x13 26      ====        srai s0, a3, 26
                                                  30'd    9100    : data = 32'h    C56D0693    ;    //    addi x13 x26 -938      ====        addi a3, s10, -938
                                                  30'd    9101    : data = 32'h    01A6C633    ;    //    xor x12 x13 x26      ====        xor a2, a3, s10
                                                  30'd    9102    : data = 32'h    016218B3    ;    //    sll x17 x4 x22      ====        sll a7, tp, s6
                                                  30'd    9103    : data = 32'h    5AEAEE13    ;    //    ori x28 x21 1454      ====        ori t3, s5, 1454
                                                  30'd    9104    : data = 32'h    01D43B33    ;    //    sltu x22 x8 x29      ====        sltu s6, s0, t4
                                                  30'd    9105    : data = 32'h    41C888B3    ;    //    sub x17 x17 x28      ====        sub a7, a7, t3
                                                  30'd    9106    : data = 32'h    404A8BB3    ;    //    sub x23 x21 x4      ====        sub s7, s5, tp
                                                  30'd    9107    : data = 32'h    113A2613    ;    //    slti x12 x20 275      ====        slti a2, s4, 275
                                                  30'd    9108    : data = 32'h    005B5833    ;    //    srl x16 x22 x5      ====        srl a6, s6, t0
                                                  30'd    9109    : data = 32'h    009ED293    ;    //    srli x5 x29 9      ====        srli t0, t4, 9
                                                  30'd    9110    : data = 32'h    3263B113    ;    //    sltiu x2 x7 806      ====        sltiu sp, t2, 806
                                                  30'd    9111    : data = 32'h    015809B3    ;    //    add x19 x16 x21      ====        add s3, a6, s5
                                                  30'd    9112    : data = 32'h    E8464897    ;    //    auipc x17 951396      ====        auipc a7, 951396
                                                  30'd    9113    : data = 32'h    3A32AF93    ;    //    slti x31 x5 931      ====        slti t6, t0, 931
                                                  30'd    9114    : data = 32'h    ED8E2393    ;    //    slti x7 x28 -296      ====        slti t2, t3, -296
                                                  30'd    9115    : data = 32'h    0062BFB3    ;    //    sltu x31 x5 x6      ====        sltu t6, t0, t1
                                                  30'd    9116    : data = 32'h    003B6933    ;    //    or x18 x22 x3      ====        or s2, s6, gp
                                                  30'd    9117    : data = 32'h    0081A033    ;    //    slt x0 x3 x8      ====        slt zero, gp, s0
                                                  30'd    9118    : data = 32'h    B3B64E13    ;    //    xori x28 x12 -1221      ====        xori t3, a2, -1221
                                                  30'd    9119    : data = 32'h    00771E13    ;    //    slli x28 x14 7      ====        slli t3, a4, 7
                                                  30'd    9120    : data = 32'h    00F0E4B3    ;    //    or x9 x1 x15      ====        or s1, ra, a5
                                                  30'd    9121    : data = 32'h    00CC76B3    ;    //    and x13 x24 x12      ====        and a3, s8, a2
                                                  30'd    9122    : data = 32'h    431D6013    ;    //    ori x0 x26 1073      ====        ori zero, s10, 1073
                                                  30'd    9123    : data = 32'h    20760813    ;    //    addi x16 x12 519      ====        addi a6, a2, 519
                                                  30'd    9124    : data = 32'h    19EDE913    ;    //    ori x18 x27 414      ====        ori s2, s11, 414
                                                  30'd    9125    : data = 32'h    5FE44637    ;    //    lui x12 392772      ====        lui a2, 392772
                                                  30'd    9126    : data = 32'h    00535C13    ;    //    srli x24 x6 5      ====        srli s8, t1, 5
                                                  30'd    9127    : data = 32'h    01E086B3    ;    //    add x13 x1 x30      ====        add a3, ra, t5
                                                  30'd    9128    : data = 32'h    9FAA4293    ;    //    xori x5 x20 -1542      ====        xori t0, s4, -1542
                                                  30'd    9129    : data = 32'h    4021D493    ;    //    srai x9 x3 2      ====        srai s1, gp, 2
                                                  30'd    9130    : data = 32'h    8B726A13    ;    //    ori x20 x4 -1865      ====        ori s4, tp, -1865
                                                  30'd    9131    : data = 32'h    019818B3    ;    //    sll x17 x16 x25      ====        sll a7, a6, s9
                                                  30'd    9132    : data = 32'h    01D641B3    ;    //    xor x3 x12 x29      ====        xor gp, a2, t4
                                                  30'd    9133    : data = 32'h    41C55893    ;    //    srai x17 x10 28      ====        srai a7, a0, 28
                                                  30'd    9134    : data = 32'h    8723EC13    ;    //    ori x24 x7 -1934      ====        ori s8, t2, -1934
                                                  30'd    9135    : data = 32'h    3BF9E593    ;    //    ori x11 x19 959      ====        ori a1, s3, 959
                                                  30'd    9136    : data = 32'h    401EDE93    ;    //    srai x29 x29 1      ====        srai t4, t4, 1
                                                  30'd    9137    : data = 32'h    CA2C0D13    ;    //    addi x26 x24 -862      ====        addi s10, s8, -862
                                                  30'd    9138    : data = 32'h    414A80B3    ;    //    sub x1 x21 x20      ====        sub ra, s5, s4
                                                  30'd    9139    : data = 32'h    401AD413    ;    //    srai x8 x21 1      ====        srai s0, s5, 1
                                                  30'd    9140    : data = 32'h    8F97A893    ;    //    slti x17 x15 -1799      ====        slti a7, a5, -1799
                                                  30'd    9141    : data = 32'h    AF814693    ;    //    xori x13 x2 -1288      ====        xori a3, sp, -1288
                                                  30'd    9142    : data = 32'h    01028E33    ;    //    add x28 x5 x16      ====        add t3, t0, a6
                                                  30'd    9143    : data = 32'h    4891CE93    ;    //    xori x29 x3 1161      ====        xori t4, gp, 1161
                                                  30'd    9144    : data = 32'h    E645A713    ;    //    slti x14 x11 -412      ====        slti a4, a1, -412
                                                  30'd    9145    : data = 32'h    65AB4993    ;    //    xori x19 x22 1626      ====        xori s3, s6, 1626
                                                  30'd    9146    : data = 32'h    6A1B7813    ;    //    andi x16 x22 1697      ====        andi a6, s6, 1697
                                                  30'd    9147    : data = 32'h    01D37733    ;    //    and x14 x6 x29      ====        and a4, t1, t4
                                                  30'd    9148    : data = 32'h    4A91A693    ;    //    slti x13 x3 1193      ====        slti a3, gp, 1193
                                                  30'd    9149    : data = 32'h    41C90FB3    ;    //    sub x31 x18 x28      ====        sub t6, s2, t3
                                                  30'd    9150    : data = 32'h    017D77B3    ;    //    and x15 x26 x23      ====        and a5, s10, s7
                                                  30'd    9151    : data = 32'h    01445893    ;    //    srli x17 x8 20      ====        srli a7, s0, 20
                                                  30'd    9152    : data = 32'h    00F41B33    ;    //    sll x22 x8 x15      ====        sll s6, s0, a5
                                                  30'd    9153    : data = 32'h    01D7A4B3    ;    //    slt x9 x15 x29      ====        slt s1, a5, t4
                                                  30'd    9154    : data = 32'h    01306633    ;    //    or x12 x0 x19      ====        or a2, zero, s3
                                                  30'd    9155    : data = 32'h    A04BA093    ;    //    slti x1 x23 -1532      ====        slti ra, s7, -1532
                                                  30'd    9156    : data = 32'h    19B18A13    ;    //    addi x20 x3 411      ====        addi s4, gp, 411
                                                  30'd    9157    : data = 32'h    E2727317    ;    //    auipc x6 927527      ====        auipc t1, 927527
                                                  30'd    9158    : data = 32'h    016BBFB3    ;    //    sltu x31 x23 x22      ====        sltu t6, s7, s6
                                                  30'd    9159    : data = 32'h    BF31BB93    ;    //    sltiu x23 x3 -1037      ====        sltiu s7, gp, -1037
                                                  30'd    9160    : data = 32'h    A1C9F893    ;    //    andi x17 x19 -1508      ====        andi a7, s3, -1508
                                                  30'd    9161    : data = 32'h    5EFEE913    ;    //    ori x18 x29 1519      ====        ori s2, t4, 1519
                                                  30'd    9162    : data = 32'h    01EE37B3    ;    //    sltu x15 x28 x30      ====        sltu a5, t3, t5
                                                  30'd    9163    : data = 32'h    CC4F3093    ;    //    sltiu x1 x30 -828      ====        sltiu ra, t5, -828
                                                  30'd    9164    : data = 32'h    13CC4613    ;    //    xori x12 x24 316      ====        xori a2, s8, 316
                                                  30'd    9165    : data = 32'h    A3D8FC93    ;    //    andi x25 x17 -1475      ====        andi s9, a7, -1475
                                                  30'd    9166    : data = 32'h    5360F393    ;    //    andi x7 x1 1334      ====        andi t2, ra, 1334
                                                  30'd    9167    : data = 32'h    000E57B3    ;    //    srl x15 x28 x0      ====        srl a5, t3, zero
                                                  30'd    9168    : data = 32'h    41EC82B3    ;    //    sub x5 x25 x30      ====        sub t0, s9, t5
                                                  30'd    9169    : data = 32'h    40AB5933    ;    //    sra x18 x22 x10      ====        sra s2, s6, a0
                                                  30'd    9170    : data = 32'h    411AEE13    ;    //    ori x28 x21 1041      ====        ori t3, s5, 1041
                                                  30'd    9171    : data = 32'h    01897CB3    ;    //    and x25 x18 x24      ====        and s9, s2, s8
                                                  30'd    9172    : data = 32'h    010E9633    ;    //    sll x12 x29 x16      ====        sll a2, t4, a6
                                                  30'd    9173    : data = 32'h    010BE633    ;    //    or x12 x23 x16      ====        or a2, s7, a6
                                                  30'd    9174    : data = 32'h    41F853B3    ;    //    sra x7 x16 x31      ====        sra t2, a6, t6
                                                  30'd    9175    : data = 32'h    DBF62A93    ;    //    slti x21 x12 -577      ====        slti s5, a2, -577
                                                  30'd    9176    : data = 32'h    01373EB3    ;    //    sltu x29 x14 x19      ====        sltu t4, a4, s3
                                                  30'd    9177    : data = 32'h    1BC2E593    ;    //    ori x11 x5 444      ====        ori a1, t0, 444
                                                  30'd    9178    : data = 32'h    01119C93    ;    //    slli x25 x3 17      ====        slli s9, gp, 17
                                                  30'd    9179    : data = 32'h    001201B3    ;    //    add x3 x4 x1      ====        add gp, tp, ra
                                                  30'd    9180    : data = 32'h    8B794793    ;    //    xori x15 x18 -1865      ====        xori a5, s2, -1865
                                                  30'd    9181    : data = 32'h    418A54B3    ;    //    sra x9 x20 x24      ====        sra s1, s4, s8
                                                  30'd    9182    : data = 32'h    00E1E1B3    ;    //    or x3 x3 x14      ====        or gp, gp, a4
                                                  30'd    9183    : data = 32'h    402C8833    ;    //    sub x16 x25 x2      ====        sub a6, s9, sp
                                                  30'd    9184    : data = 32'h    B35D0113    ;    //    addi x2 x26 -1227      ====        addi sp, s10, -1227
                                                  30'd    9185    : data = 32'h    008D5913    ;    //    srli x18 x26 8      ====        srli s2, s10, 8
                                                  30'd    9186    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9187    : data = 32'h    D55F3993    ;    //    sltiu x19 x30 -683      ====        sltiu s3, t5, -683
                                                  30'd    9188    : data = 32'h    3BF67B17    ;    //    auipc x22 245607      ====        auipc s6, 245607
                                                  30'd    9189    : data = 32'h    011A83B3    ;    //    add x7 x21 x17      ====        add t2, s5, a7
                                                  30'd    9190    : data = 32'h    40D4D9B3    ;    //    sra x19 x9 x13      ====        sra s3, s1, a3
                                                  30'd    9191    : data = 32'h    5B7B6E13    ;    //    ori x28 x22 1463      ====        ori t3, s6, 1463
                                                  30'd    9192    : data = 32'h    01A8B4B3    ;    //    sltu x9 x17 x26      ====        sltu s1, a7, s10
                                                  30'd    9193    : data = 32'h    CF1AB713    ;    //    sltiu x14 x21 -783      ====        sltiu a4, s5, -783
                                                  30'd    9194    : data = 32'h    A06D6B93    ;    //    ori x23 x26 -1530      ====        ori s7, s10, -1530
                                                  30'd    9195    : data = 32'h    DB31BD93    ;    //    sltiu x27 x3 -589      ====        sltiu s11, gp, -589
                                                  30'd    9196    : data = 32'h    6797CB13    ;    //    xori x22 x15 1657      ====        xori s6, a5, 1657
                                                  30'd    9197    : data = 32'h    00E06333    ;    //    or x6 x0 x14      ====        or t1, zero, a4
                                                  30'd    9198    : data = 32'h    22E8C393    ;    //    xori x7 x17 558      ====        xori t2, a7, 558
                                                  30'd    9199    : data = 32'h    019F1E93    ;    //    slli x29 x30 25      ====        slli t4, t5, 25
                                                  30'd    9200    : data = 32'h    0186F633    ;    //    and x12 x13 x24      ====        and a2, a3, s8
                                                  30'd    9201    : data = 32'h    645CBE13    ;    //    sltiu x28 x25 1605      ====        sltiu t3, s9, 1605
                                                  30'd    9202    : data = 32'h    D6060313    ;    //    addi x6 x12 -672      ====        addi t1, a2, -672
                                                  30'd    9203    : data = 32'h    40B55613    ;    //    srai x12 x10 11      ====        srai a2, a0, 11
                                                  30'd    9204    : data = 32'h    00144D33    ;    //    xor x26 x8 x1      ====        xor s10, s0, ra
                                                  30'd    9205    : data = 32'h    41E7DBB3    ;    //    sra x23 x15 x30      ====        sra s7, a5, t5
                                                  30'd    9206    : data = 32'h    B74B7B13    ;    //    andi x22 x22 -1164      ====        andi s6, s6, -1164
                                                  30'd    9207    : data = 32'h    54630F93    ;    //    addi x31 x6 1350      ====        addi t6, t1, 1350
                                                  30'd    9208    : data = 32'h    414E0633    ;    //    sub x12 x28 x20      ====        sub a2, t3, s4
                                                  30'd    9209    : data = 32'h    CD53A2B7    ;    //    lui x5 841018      ====        lui t0, 841018
                                                  30'd    9210    : data = 32'h    41A05D13    ;    //    srai x26 x0 26      ====        srai s10, zero, 26
                                                  30'd    9211    : data = 32'h    004A8933    ;    //    add x18 x21 x4      ====        add s2, s5, tp
                                                  30'd    9212    : data = 32'h    C9F14993    ;    //    xori x19 x2 -865      ====        xori s3, sp, -865
                                                  30'd    9213    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9214    : data = 32'h    30F83713    ;    //    sltiu x14 x16 783      ====        sltiu a4, a6, 783
                                                  30'd    9215    : data = 32'h    F5D1D297    ;    //    auipc x5 1006877      ====        auipc t0, 1006877
                                                  30'd    9216    : data = 32'h    49648713    ;    //    addi x14 x9 1174      ====        addi a4, s1, 1174
                                                  30'd    9217    : data = 32'h    27BAE393    ;    //    ori x7 x21 635      ====        ori t2, s5, 635
                                                  30'd    9218    : data = 32'h    01257933    ;    //    and x18 x10 x18      ====        and s2, a0, s2
                                                  30'd    9219    : data = 32'h    0740B893    ;    //    sltiu x17 x1 116      ====        sltiu a7, ra, 116
                                                  30'd    9220    : data = 32'h    24BBEA17    ;    //    auipc x20 150462      ====        auipc s4, 150462
                                                  30'd    9221    : data = 32'h    4571F997    ;    //    auipc x19 284447      ====        auipc s3, 284447
                                                  30'd    9222    : data = 32'h    01CAF5B3    ;    //    and x11 x21 x28      ====        and a1, s5, t3
                                                  30'd    9223    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9224    : data = 32'h    2479CE13    ;    //    xori x28 x19 583      ====        xori t3, s3, 583
                                                  30'd    9225    : data = 32'h    01C3D633    ;    //    srl x12 x7 x28      ====        srl a2, t2, t3
                                                  30'd    9226    : data = 32'h    42540793    ;    //    addi x15 x8 1061      ====        addi a5, s0, 1061
                                                  30'd    9227    : data = 32'h    01C611B3    ;    //    sll x3 x12 x28      ====        sll gp, a2, t3
                                                  30'd    9228    : data = 32'h    3D73A813    ;    //    slti x16 x7 983      ====        slti a6, t2, 983
                                                  30'd    9229    : data = 32'h    BD951697    ;    //    auipc x13 776529      ====        auipc a3, 776529
                                                  30'd    9230    : data = 32'h    670AFA13    ;    //    andi x20 x21 1648      ====        andi s4, s5, 1648
                                                  30'd    9231    : data = 32'h    40375AB3    ;    //    sra x21 x14 x3      ====        sra s5, a4, gp
                                                  30'd    9232    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9233    : data = 32'h    0126E633    ;    //    or x12 x13 x18      ====        or a2, a3, s2
                                                  30'd    9234    : data = 32'h    01B3E1B3    ;    //    or x3 x7 x27      ====        or gp, t2, s11
                                                  30'd    9235    : data = 32'h    003ED133    ;    //    srl x2 x29 x3      ====        srl sp, t4, gp
                                                  30'd    9236    : data = 32'h    41DD5F93    ;    //    srai x31 x26 29      ====        srai t6, s10, 29
                                                  30'd    9237    : data = 32'h    F44CE113    ;    //    ori x2 x25 -188      ====        ori sp, s9, -188
                                                  30'd    9238    : data = 32'h    01D24E33    ;    //    xor x28 x4 x29      ====        xor t3, tp, t4
                                                  30'd    9239    : data = 32'h    41DA5833    ;    //    sra x16 x20 x29      ====        sra a6, s4, t4
                                                  30'd    9240    : data = 32'h    7BB298B7    ;    //    lui x17 506665      ====        lui a7, 506665
                                                  30'd    9241    : data = 32'h    01649133    ;    //    sll x2 x9 x22      ====        sll sp, s1, s6
                                                  30'd    9242    : data = 32'h    00A13433    ;    //    sltu x8 x2 x10      ====        sltu s0, sp, a0
                                                  30'd    9243    : data = 32'h    EF4DFF93    ;    //    andi x31 x27 -268      ====        andi t6, s11, -268
                                                  30'd    9244    : data = 32'h    018ED813    ;    //    srli x16 x29 24      ====        srli a6, t4, 24
                                                  30'd    9245    : data = 32'h    AD019597    ;    //    auipc x11 708633      ====        auipc a1, 708633
                                                  30'd    9246    : data = 32'h    00ED1293    ;    //    slli x5 x26 14      ====        slli t0, s10, 14
                                                  30'd    9247    : data = 32'h    012C0D33    ;    //    add x26 x24 x18      ====        add s10, s8, s2
                                                  30'd    9248    : data = 32'h    000344B3    ;    //    xor x9 x6 x0      ====        xor s1, t1, zero
                                                  30'd    9249    : data = 32'h    0178ECB3    ;    //    or x25 x17 x23      ====        or s9, a7, s7
                                                  30'd    9250    : data = 32'h    00B91693    ;    //    slli x13 x18 11      ====        slli a3, s2, 11
                                                  30'd    9251    : data = 32'h    01F99A33    ;    //    sll x20 x19 x31      ====        sll s4, s3, t6
                                                  30'd    9252    : data = 32'h    DE7BDFB7    ;    //    lui x31 911293      ====        lui t6, 911293
                                                  30'd    9253    : data = 32'h    1BD4B093    ;    //    sltiu x1 x9 445      ====        sltiu ra, s1, 445
                                                  30'd    9254    : data = 32'h    0056D4B3    ;    //    srl x9 x13 x5      ====        srl s1, a3, t0
                                                  30'd    9255    : data = 32'h    AFF54613    ;    //    xori x12 x10 -1281      ====        xori a2, a0, -1281
                                                  30'd    9256    : data = 32'h    0128AD33    ;    //    slt x26 x17 x18      ====        slt s10, a7, s2
                                                  30'd    9257    : data = 32'h    D3823813    ;    //    sltiu x16 x4 -712      ====        sltiu a6, tp, -712
                                                  30'd    9258    : data = 32'h    4045D713    ;    //    srai x14 x11 4      ====        srai a4, a1, 4
                                                  30'd    9259    : data = 32'h    0181BB33    ;    //    sltu x22 x3 x24      ====        sltu s6, gp, s8
                                                  30'd    9260    : data = 32'h    40D75D13    ;    //    srai x26 x14 13      ====        srai s10, a4, 13
                                                  30'd    9261    : data = 32'h    018AFCB3    ;    //    and x25 x21 x24      ====        and s9, s5, s8
                                                  30'd    9262    : data = 32'h    40560633    ;    //    sub x12 x12 x5      ====        sub a2, a2, t0
                                                  30'd    9263    : data = 32'h    01284633    ;    //    xor x12 x16 x18      ====        xor a2, a6, s2
                                                  30'd    9264    : data = 32'h    00BE3733    ;    //    sltu x14 x28 x11      ====        sltu a4, t3, a1
                                                  30'd    9265    : data = 32'h    002E9133    ;    //    sll x2 x29 x2      ====        sll sp, t4, sp
                                                  30'd    9266    : data = 32'h    00031393    ;    //    slli x7 x6 0      ====        slli t2, t1, 0
                                                  30'd    9267    : data = 32'h    017EDA13    ;    //    srli x20 x29 23      ====        srli s4, t4, 23
                                                  30'd    9268    : data = 32'h    00C39C93    ;    //    slli x25 x7 12      ====        slli s9, t2, 12
                                                  30'd    9269    : data = 32'h    00A589B3    ;    //    add x19 x11 x10      ====        add s3, a1, a0
                                                  30'd    9270    : data = 32'h    01423FB3    ;    //    sltu x31 x4 x20      ====        sltu t6, tp, s4
                                                  30'd    9271    : data = 32'h    013C79B3    ;    //    and x19 x24 x19      ====        and s3, s8, s3
                                                  30'd    9272    : data = 32'h    011FEFB3    ;    //    or x31 x31 x17      ====        or t6, t6, a7
                                                  30'd    9273    : data = 32'h    01A7AEB3    ;    //    slt x29 x15 x26      ====        slt t4, a5, s10
                                                  30'd    9274    : data = 32'h    014DC9B3    ;    //    xor x19 x27 x20      ====        xor s3, s11, s4
                                                  30'd    9275    : data = 32'h    1C256097    ;    //    auipc x1 115286      ====        auipc ra, 115286
                                                  30'd    9276    : data = 32'h    01884833    ;    //    xor x16 x16 x24      ====        xor a6, a6, s8
                                                  30'd    9277    : data = 32'h    00893E33    ;    //    sltu x28 x18 x8      ====        sltu t3, s2, s0
                                                  30'd    9278    : data = 32'h    01D3BC33    ;    //    sltu x24 x7 x29      ====        sltu s8, t2, t4
                                                  30'd    9279    : data = 32'h    00DA91B3    ;    //    sll x3 x21 x13      ====        sll gp, s5, a3
                                                  30'd    9280    : data = 32'h    00B972B3    ;    //    and x5 x18 x11      ====        and t0, s2, a1
                                                  30'd    9281    : data = 32'h    DE346A97    ;    //    auipc x21 910150      ====        auipc s5, 910150
                                                  30'd    9282    : data = 32'h    010E3B33    ;    //    sltu x22 x28 x16      ====        sltu s6, t3, a6
                                                  30'd    9283    : data = 32'h    85103593    ;    //    sltiu x11 x0 -1967      ====        sltiu a1, zero, -1967
                                                  30'd    9284    : data = 32'h    00A31113    ;    //    slli x2 x6 10      ====        slli sp, t1, 10
                                                  30'd    9285    : data = 32'h    00A728B3    ;    //    slt x17 x14 x10      ====        slt a7, a4, a0
                                                  30'd    9286    : data = 32'h    6F26F593    ;    //    andi x11 x13 1778      ====        andi a1, a3, 1778
                                                  30'd    9287    : data = 32'h    00B474B3    ;    //    and x9 x8 x11      ====        and s1, s0, a1
                                                  30'd    9288    : data = 32'h    3765F613    ;    //    andi x12 x11 886      ====        andi a2, a1, 886
                                                  30'd    9289    : data = 32'h    5408E693    ;    //    ori x13 x17 1344      ====        ori a3, a7, 1344
                                                  30'd    9290    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9291    : data = 32'h    01151E93    ;    //    slli x29 x10 17      ====        slli t4, a0, 17
                                                  30'd    9292    : data = 32'h    9D0AFC93    ;    //    andi x25 x21 -1584      ====        andi s9, s5, -1584
                                                  30'd    9293    : data = 32'h    00AA2DB3    ;    //    slt x27 x20 x10      ====        slt s11, s4, a0
                                                  30'd    9294    : data = 32'h    010B75B3    ;    //    and x11 x22 x16      ====        and a1, s6, a6
                                                  30'd    9295    : data = 32'h    00956BB3    ;    //    or x23 x10 x9      ====        or s7, a0, s1
                                                  30'd    9296    : data = 32'h    40E95FB3    ;    //    sra x31 x18 x14      ====        sra t6, s2, a4
                                                  30'd    9297    : data = 32'h    01071133    ;    //    sll x2 x14 x16      ====        sll sp, a4, a6
                                                  30'd    9298    : data = 32'h    0151A033    ;    //    slt x0 x3 x21      ====        slt zero, gp, s5
                                                  30'd    9299    : data = 32'h    41360833    ;    //    sub x16 x12 x19      ====        sub a6, a2, s3
                                                  30'd    9300    : data = 32'h    41F85013    ;    //    srai x0 x16 31      ====        srai zero, a6, 31
                                                  30'd    9301    : data = 32'h    41CF5B33    ;    //    sra x22 x30 x28      ====        sra s6, t5, t3
                                                  30'd    9302    : data = 32'h    01667833    ;    //    and x16 x12 x22      ====        and a6, a2, s6
                                                  30'd    9303    : data = 32'h    75718313    ;    //    addi x6 x3 1879      ====        addi t1, gp, 1879
                                                  30'd    9304    : data = 32'h    403700B3    ;    //    sub x1 x14 x3      ====        sub ra, a4, gp
                                                  30'd    9305    : data = 32'h    4058F013    ;    //    andi x0 x17 1029      ====        andi zero, a7, 1029
                                                  30'd    9306    : data = 32'h    01E3DB33    ;    //    srl x22 x7 x30      ====        srl s6, t2, t5
                                                  30'd    9307    : data = 32'h    00FAD193    ;    //    srli x3 x21 15      ====        srli gp, s5, 15
                                                  30'd    9308    : data = 32'h    0012FD33    ;    //    and x26 x5 x1      ====        and s10, t0, ra
                                                  30'd    9309    : data = 32'h    48090E97    ;    //    auipc x29 295056      ====        auipc t4, 295056
                                                  30'd    9310    : data = 32'h    9ADBA293    ;    //    slti x5 x23 -1619      ====        slti t0, s7, -1619
                                                  30'd    9311    : data = 32'h    41290933    ;    //    sub x18 x18 x18      ====        sub s2, s2, s2
                                                  30'd    9312    : data = 32'h    004322B3    ;    //    slt x5 x6 x4      ====        slt t0, t1, tp
                                                  30'd    9313    : data = 32'h    012DBBB3    ;    //    sltu x23 x27 x18      ====        sltu s7, s11, s2
                                                  30'd    9314    : data = 32'h    F90BBD13    ;    //    sltiu x26 x23 -112      ====        sltiu s10, s7, -112
                                                  30'd    9315    : data = 32'h    00A73D33    ;    //    sltu x26 x14 x10      ====        sltu s10, a4, a0
                                                  30'd    9316    : data = 32'h    AC4BE313    ;    //    ori x6 x23 -1340      ====        ori t1, s7, -1340
                                                  30'd    9317    : data = 32'h    4037D2B3    ;    //    sra x5 x15 x3      ====        sra t0, a5, gp
                                                  30'd    9318    : data = 32'h    41F25313    ;    //    srai x6 x4 31      ====        srai t1, tp, 31
                                                  30'd    9319    : data = 32'h    40D18333    ;    //    sub x6 x3 x13      ====        sub t1, gp, a3
                                                  30'd    9320    : data = 32'h    018E7FB3    ;    //    and x31 x28 x24      ====        and t6, t3, s8
                                                  30'd    9321    : data = 32'h    41F45333    ;    //    sra x6 x8 x31      ====        sra t1, s0, t6
                                                  30'd    9322    : data = 32'h    41305FB3    ;    //    sra x31 x0 x19      ====        sra t6, zero, s3
                                                  30'd    9323    : data = 32'h    23566897    ;    //    auipc x17 144742      ====        auipc a7, 144742
                                                  30'd    9324    : data = 32'h    41645033    ;    //    sra x0 x8 x22      ====        sra zero, s0, s6
                                                  30'd    9325    : data = 32'h    012993B3    ;    //    sll x7 x19 x18      ====        sll t2, s3, s2
                                                  30'd    9326    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9327    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9328    : data = 32'h    018ED733    ;    //    srl x14 x29 x24      ====        srl a4, t4, s8
                                                  30'd    9329    : data = 32'h    01E48B33    ;    //    add x22 x9 x30      ====        add s6, s1, t5
                                                  30'd    9330    : data = 32'h    0093C3B3    ;    //    xor x7 x7 x9      ====        xor t2, t2, s1
                                                  30'd    9331    : data = 32'h    403E5293    ;    //    srai x5 x28 3      ====        srai t0, t3, 3
                                                  30'd    9332    : data = 32'h    005A9633    ;    //    sll x12 x21 x5      ====        sll a2, s5, t0
                                                  30'd    9333    : data = 32'h    77BAE893    ;    //    ori x17 x21 1915      ====        ori a7, s5, 1915
                                                  30'd    9334    : data = 32'h    415CD1B3    ;    //    sra x3 x25 x21      ====        sra gp, s9, s5
                                                  30'd    9335    : data = 32'h    414B0EB3    ;    //    sub x29 x22 x20      ====        sub t4, s6, s4
                                                  30'd    9336    : data = 32'h    2AED6717    ;    //    auipc x14 175830      ====        auipc a4, 175830
                                                  30'd    9337    : data = 32'h    E7C7C393    ;    //    xori x7 x15 -388      ====        xori t2, a5, -388
                                                  30'd    9338    : data = 32'h    41B05C33    ;    //    sra x24 x0 x27      ====        sra s8, zero, s11
                                                  30'd    9339    : data = 32'h    66203893    ;    //    sltiu x17 x0 1634      ====        sltiu a7, zero, 1634
                                                  30'd    9340    : data = 32'h    016D9A33    ;    //    sll x20 x27 x22      ====        sll s4, s11, s6
                                                  30'd    9341    : data = 32'h    019C6833    ;    //    or x16 x24 x25      ====        or a6, s8, s9
                                                  30'd    9342    : data = 32'h    FAD62113    ;    //    slti x2 x12 -83      ====        slti sp, a2, -83
                                                  30'd    9343    : data = 32'h    01952633    ;    //    slt x12 x10 x25      ====        slt a2, a0, s9
                                                  30'd    9344    : data = 32'h    00A0D113    ;    //    srli x2 x1 10      ====        srli sp, ra, 10
                                                  30'd    9345    : data = 32'h    417E5193    ;    //    srai x3 x28 23      ====        srai gp, t3, 23
                                                  30'd    9346    : data = 32'h    41FE8993    ;    //    addi x19 x29 1055      ====        addi s3, t4, 1055
                                                  30'd    9347    : data = 32'h    B19D8F93    ;    //    addi x31 x27 -1255      ====        addi t6, s11, -1255
                                                  30'd    9348    : data = 32'h    00661313    ;    //    slli x6 x12 6      ====        slli t1, a2, 6
                                                  30'd    9349    : data = 32'h    2BEAF493    ;    //    andi x9 x21 702      ====        andi s1, s5, 702
                                                  30'd    9350    : data = 32'h    002E96B3    ;    //    sll x13 x29 x2      ====        sll a3, t4, sp
                                                  30'd    9351    : data = 32'h    01F67CB3    ;    //    and x25 x12 x31      ====        and s9, a2, t6
                                                  30'd    9352    : data = 32'h    5D95FD13    ;    //    andi x26 x11 1497      ====        andi s10, a1, 1497
                                                  30'd    9353    : data = 32'h    BE1BB593    ;    //    sltiu x11 x23 -1055      ====        sltiu a1, s7, -1055
                                                  30'd    9354    : data = 32'h    A6D5AE13    ;    //    slti x28 x11 -1427      ====        slti t3, a1, -1427
                                                  30'd    9355    : data = 32'h    905BA637    ;    //    lui x12 591290      ====        lui a2, 591290
                                                  30'd    9356    : data = 32'h    41E8D633    ;    //    sra x12 x17 x30      ====        sra a2, a7, t5
                                                  30'd    9357    : data = 32'h    CCB16B17    ;    //    auipc x22 838422      ====        auipc s6, 838422
                                                  30'd    9358    : data = 32'h    1D1DF313    ;    //    andi x6 x27 465      ====        andi t1, s11, 465
                                                  30'd    9359    : data = 32'h    38F9C793    ;    //    xori x15 x19 911      ====        xori a5, s3, 911
                                                  30'd    9360    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9361    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9362    : data = 32'h    012EAAB3    ;    //    slt x21 x29 x18      ====        slt s5, t4, s2
                                                  30'd    9363    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9364    : data = 32'h    00F220B3    ;    //    slt x1 x4 x15      ====        slt ra, tp, a5
                                                  30'd    9365    : data = 32'h    01279393    ;    //    slli x7 x15 18      ====        slli t2, a5, 18
                                                  30'd    9366    : data = 32'h    009023B3    ;    //    slt x7 x0 x9      ====        slt t2, zero, s1
                                                  30'd    9367    : data = 32'h    0175EE33    ;    //    or x28 x11 x23      ====        or t3, a1, s7
                                                  30'd    9368    : data = 32'h    9575C313    ;    //    xori x6 x11 -1705      ====        xori t1, a1, -1705
                                                  30'd    9369    : data = 32'h    405AD713    ;    //    srai x14 x21 5      ====        srai a4, s5, 5
                                                  30'd    9370    : data = 32'h    0136E7B3    ;    //    or x15 x13 x19      ====        or a5, a3, s3
                                                  30'd    9371    : data = 32'h    00661313    ;    //    slli x6 x12 6      ====        slli t1, a2, 6
                                                  30'd    9372    : data = 32'h    0148D4B3    ;    //    srl x9 x17 x20      ====        srl s1, a7, s4
                                                  30'd    9373    : data = 32'h    0178D693    ;    //    srli x13 x17 23      ====        srli a3, a7, 23
                                                  30'd    9374    : data = 32'h    00D10133    ;    //    add x2 x2 x13      ====        add sp, sp, a3
                                                  30'd    9375    : data = 32'h    0057C9B3    ;    //    xor x19 x15 x5      ====        xor s3, a5, t0
                                                  30'd    9376    : data = 32'h    40145713    ;    //    srai x14 x8 1      ====        srai a4, s0, 1
                                                  30'd    9377    : data = 32'h    005DE833    ;    //    or x16 x27 x5      ====        or a6, s11, t0
                                                  30'd    9378    : data = 32'h    E2A7C413    ;    //    xori x8 x15 -470      ====        xori s0, a5, -470
                                                  30'd    9379    : data = 32'h    01977FB3    ;    //    and x31 x14 x25      ====        and t6, a4, s9
                                                  30'd    9380    : data = 32'h    0D739F97    ;    //    auipc x31 55097      ====        auipc t6, 55097
                                                  30'd    9381    : data = 32'h    D4622C13    ;    //    slti x24 x4 -698      ====        slti s8, tp, -698
                                                  30'd    9382    : data = 32'h    01EDDD13    ;    //    srli x26 x27 30      ====        srli s10, s11, 30
                                                  30'd    9383    : data = 32'h    40975EB3    ;    //    sra x29 x14 x9      ====        sra t4, a4, s1
                                                  30'd    9384    : data = 32'h    00387333    ;    //    and x6 x16 x3      ====        and t1, a6, gp
                                                  30'd    9385    : data = 32'h    2284B193    ;    //    sltiu x3 x9 552      ====        sltiu gp, s1, 552
                                                  30'd    9386    : data = 32'h    892BAD13    ;    //    slti x26 x23 -1902      ====        slti s10, s7, -1902
                                                  30'd    9387    : data = 32'h    F66C6393    ;    //    ori x7 x24 -154      ====        ori t2, s8, -154
                                                  30'd    9388    : data = 32'h    41D80BB3    ;    //    sub x23 x16 x29      ====        sub s7, a6, t4
                                                  30'd    9389    : data = 32'h    01B44433    ;    //    xor x8 x8 x27      ====        xor s0, s0, s11
                                                  30'd    9390    : data = 32'h    40910CB3    ;    //    sub x25 x2 x9      ====        sub s9, sp, s1
                                                  30'd    9391    : data = 32'h    00D519B3    ;    //    sll x19 x10 x13      ====        sll s3, a0, a3
                                                  30'd    9392    : data = 32'h    7964FB13    ;    //    andi x22 x9 1942      ====        andi s6, s1, 1942
                                                  30'd    9393    : data = 32'h    27FDC613    ;    //    xori x12 x27 639      ====        xori a2, s11, 639
                                                  30'd    9394    : data = 32'h    8F58FC93    ;    //    andi x25 x17 -1803      ====        andi s9, a7, -1803
                                                  30'd    9395    : data = 32'h    01E41D33    ;    //    sll x26 x8 x30      ====        sll s10, s0, t5
                                                  30'd    9396    : data = 32'h    40A35433    ;    //    sra x8 x6 x10      ====        sra s0, t1, a0
                                                  30'd    9397    : data = 32'h    01239A13    ;    //    slli x20 x7 18      ====        slli s4, t2, 18
                                                  30'd    9398    : data = 32'h    4167D033    ;    //    sra x0 x15 x22      ====        sra zero, a5, s6
                                                  30'd    9399    : data = 32'h    F0143113    ;    //    sltiu x2 x8 -255      ====        sltiu sp, s0, -255
                                                  30'd    9400    : data = 32'h    154A4E13    ;    //    xori x28 x20 340      ====        xori t3, s4, 340
                                                  30'd    9401    : data = 32'h    014D5793    ;    //    srli x15 x26 20      ====        srli a5, s10, 20
                                                  30'd    9402    : data = 32'h    DF779BB7    ;    //    lui x23 915321      ====        lui s7, 915321
                                                  30'd    9403    : data = 32'h    01621033    ;    //    sll x0 x4 x22      ====        sll zero, tp, s6
                                                  30'd    9404    : data = 32'h    01367BB3    ;    //    and x23 x12 x19      ====        and s7, a2, s3
                                                  30'd    9405    : data = 32'h    E9A44A13    ;    //    xori x20 x8 -358      ====        xori s4, s0, -358
                                                  30'd    9406    : data = 32'h    407ED393    ;    //    srai x7 x29 7      ====        srai t2, t4, 7
                                                  30'd    9407    : data = 32'h    A00E7E13    ;    //    andi x28 x28 -1536      ====        andi t3, t3, -1536
                                                  30'd    9408    : data = 32'h    CD4FF793    ;    //    andi x15 x31 -812      ====        andi a5, t6, -812
                                                  30'd    9409    : data = 32'h    011DF3B3    ;    //    and x7 x27 x17      ====        and t2, s11, a7
                                                  30'd    9410    : data = 32'h    01552A33    ;    //    slt x20 x10 x21      ====        slt s4, a0, s5
                                                  30'd    9411    : data = 32'h    00C2FB33    ;    //    and x22 x5 x12      ====        and s6, t0, a2
                                                  30'd    9412    : data = 32'h    0C28F713    ;    //    andi x14 x17 194      ====        andi a4, a7, 194
                                                  30'd    9413    : data = 32'h    9F9D4F93    ;    //    xori x31 x26 -1543      ====        xori t6, s10, -1543
                                                  30'd    9414    : data = 32'h    019BEB33    ;    //    or x22 x23 x25      ====        or s6, s7, s9
                                                  30'd    9415    : data = 32'h    405BF1B7    ;    //    lui x3 263615      ====        lui gp, 263615
                                                  30'd    9416    : data = 32'h    40A7DC13    ;    //    srai x24 x15 10      ====        srai s8, a5, 10
                                                  30'd    9417    : data = 32'h    01CE7133    ;    //    and x2 x28 x28      ====        and sp, t3, t3
                                                  30'd    9418    : data = 32'h    02EB4913    ;    //    xori x18 x22 46      ====        xori s2, s6, 46
                                                  30'd    9419    : data = 32'h    40EE8BB3    ;    //    sub x23 x29 x14      ====        sub s7, t4, a4
                                                  30'd    9420    : data = 32'h    41BD0833    ;    //    sub x16 x26 x27      ====        sub a6, s10, s11
                                                  30'd    9421    : data = 32'h    4172D293    ;    //    srai x5 x5 23      ====        srai t0, t0, 23
                                                  30'd    9422    : data = 32'h    010A8833    ;    //    add x16 x21 x16      ====        add a6, s5, a6
                                                  30'd    9423    : data = 32'h    004EDDB3    ;    //    srl x27 x29 x4      ====        srl s11, t4, tp
                                                  30'd    9424    : data = 32'h    006EA4B3    ;    //    slt x9 x29 x6      ====        slt s1, t4, t1
                                                  30'd    9425    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9426    : data = 32'h    8AC47417    ;    //    auipc x8 568391      ====        auipc s0, 568391
                                                  30'd    9427    : data = 32'h    41C156B3    ;    //    sra x13 x2 x28      ====        sra a3, sp, t3
                                                  30'd    9428    : data = 32'h    01F65413    ;    //    srli x8 x12 31      ====        srli s0, a2, 31
                                                  30'd    9429    : data = 32'h    00EEDE93    ;    //    srli x29 x29 14      ====        srli t4, t4, 14
                                                  30'd    9430    : data = 32'h    008292B3    ;    //    sll x5 x5 x8      ====        sll t0, t0, s0
                                                  30'd    9431    : data = 32'h    8AF7FF93    ;    //    andi x31 x15 -1873      ====        andi t6, a5, -1873
                                                  30'd    9432    : data = 32'h    00861033    ;    //    sll x0 x12 x8      ====        sll zero, a2, s0
                                                  30'd    9433    : data = 32'h    B29ECD37    ;    //    lui x26 731628      ====        lui s10, 731628
                                                  30'd    9434    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9435    : data = 32'h    009284B3    ;    //    add x9 x5 x9      ====        add s1, t0, s1
                                                  30'd    9436    : data = 32'h    964C0C13    ;    //    addi x24 x24 -1692      ====        addi s8, s8, -1692
                                                  30'd    9437    : data = 32'h    00D95813    ;    //    srli x16 x18 13      ====        srli a6, s2, 13
                                                  30'd    9438    : data = 32'h    FCF07893    ;    //    andi x17 x0 -49      ====        andi a7, zero, -49
                                                  30'd    9439    : data = 32'h    000AD3B3    ;    //    srl x7 x21 x0      ====        srl t2, s5, zero
                                                  30'd    9440    : data = 32'h    008013B3    ;    //    sll x7 x0 x8      ====        sll t2, zero, s0
                                                  30'd    9441    : data = 32'h    007668B3    ;    //    or x17 x12 x7      ====        or a7, a2, t2
                                                  30'd    9442    : data = 32'h    2F470117    ;    //    auipc x2 193648      ====        auipc sp, 193648
                                                  30'd    9443    : data = 32'h    001174B3    ;    //    and x9 x2 x1      ====        and s1, sp, ra
                                                  30'd    9444    : data = 32'h    00E317B3    ;    //    sll x15 x6 x14      ====        sll a5, t1, a4
                                                  30'd    9445    : data = 32'h    5D0EE393    ;    //    ori x7 x29 1488      ====        ori t2, t4, 1488
                                                  30'd    9446    : data = 32'h    00E7F5B3    ;    //    and x11 x15 x14      ====        and a1, a5, a4
                                                  30'd    9447    : data = 32'h    8A62E293    ;    //    ori x5 x5 -1882      ====        ori t0, t0, -1882
                                                  30'd    9448    : data = 32'h    017AECB3    ;    //    or x25 x21 x23      ====        or s9, s5, s7
                                                  30'd    9449    : data = 32'h    415908B3    ;    //    sub x17 x18 x21      ====        sub a7, s2, s5
                                                  30'd    9450    : data = 32'h    8EF70113    ;    //    addi x2 x14 -1809      ====        addi sp, a4, -1809
                                                  30'd    9451    : data = 32'h    AB609AB7    ;    //    lui x21 701961      ====        lui s5, 701961
                                                  30'd    9452    : data = 32'h    01E012B3    ;    //    sll x5 x0 x30      ====        sll t0, zero, t5
                                                  30'd    9453    : data = 32'h    94833C93    ;    //    sltiu x25 x6 -1720      ====        sltiu s9, t1, -1720
                                                  30'd    9454    : data = 32'h    01185313    ;    //    srli x6 x16 17      ====        srli t1, a6, 17
                                                  30'd    9455    : data = 32'h    00FAD313    ;    //    srli x6 x21 15      ====        srli t1, s5, 15
                                                  30'd    9456    : data = 32'h    6E740013    ;    //    addi x0 x8 1767      ====        addi zero, s0, 1767
                                                  30'd    9457    : data = 32'h    010C99B3    ;    //    sll x19 x25 x16      ====        sll s3, s9, a6
                                                  30'd    9458    : data = 32'h    012878B3    ;    //    and x17 x16 x18      ====        and a7, a6, s2
                                                  30'd    9459    : data = 32'h    C618B093    ;    //    sltiu x1 x17 -927      ====        sltiu ra, a7, -927
                                                  30'd    9460    : data = 32'h    652FA037    ;    //    lui x0 414458      ====        lui zero, 414458
                                                  30'd    9461    : data = 32'h    4D326993    ;    //    ori x19 x4 1235      ====        ori s3, tp, 1235
                                                  30'd    9462    : data = 32'h    004188B3    ;    //    add x17 x3 x4      ====        add a7, gp, tp
                                                  30'd    9463    : data = 32'h    00549A13    ;    //    slli x20 x9 5      ====        slli s4, s1, 5
                                                  30'd    9464    : data = 32'h    414905B3    ;    //    sub x11 x18 x20      ====        sub a1, s2, s4
                                                  30'd    9465    : data = 32'h    016DB8B3    ;    //    sltu x17 x27 x22      ====        sltu a7, s11, s6
                                                  30'd    9466    : data = 32'h    00DDB2B3    ;    //    sltu x5 x27 x13      ====        sltu t0, s11, a3
                                                  30'd    9467    : data = 32'h    41F7D293    ;    //    srai x5 x15 31      ====        srai t0, a5, 31
                                                  30'd    9468    : data = 32'h    00981593    ;    //    slli x11 x16 9      ====        slli a1, a6, 9
                                                  30'd    9469    : data = 32'h    1276B993    ;    //    sltiu x19 x13 295      ====        sltiu s3, a3, 295
                                                  30'd    9470    : data = 32'h    00A29293    ;    //    slli x5 x5 10      ====        slli t0, t0, 10
                                                  30'd    9471    : data = 32'h    21528117    ;    //    auipc x2 136488      ====        auipc sp, 136488
                                                  30'd    9472    : data = 32'h    01FF63B3    ;    //    or x7 x30 x31      ====        or t2, t5, t6
                                                  30'd    9473    : data = 32'h    00A5AB33    ;    //    slt x22 x11 x10      ====        slt s6, a1, a0
                                                  30'd    9474    : data = 32'h    008D11B3    ;    //    sll x3 x26 x8      ====        sll gp, s10, s0
                                                  30'd    9475    : data = 32'h    015D9D33    ;    //    sll x26 x27 x21      ====        sll s10, s11, s5
                                                  30'd    9476    : data = 32'h    00FE1A13    ;    //    slli x20 x28 15      ====        slli s4, t3, 15
                                                  30'd    9477    : data = 32'h    AF247193    ;    //    andi x3 x8 -1294      ====        andi gp, s0, -1294
                                                  30'd    9478    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9479    : data = 32'h    013CA733    ;    //    slt x14 x25 x19      ====        slt a4, s9, s3
                                                  30'd    9480    : data = 32'h    4186DD33    ;    //    sra x26 x13 x24      ====        sra s10, a3, s8
                                                  30'd    9481    : data = 32'h    8D5F3693    ;    //    sltiu x13 x30 -1835      ====        sltiu a3, t5, -1835
                                                  30'd    9482    : data = 32'h    8A6CC793    ;    //    xori x15 x25 -1882      ====        xori a5, s9, -1882
                                                  30'd    9483    : data = 32'h    01572C33    ;    //    slt x24 x14 x21      ====        slt s8, a4, s5
                                                  30'd    9484    : data = 32'h    404C5713    ;    //    srai x14 x24 4      ====        srai a4, s8, 4
                                                  30'd    9485    : data = 32'h    0128F0B3    ;    //    and x1 x17 x18      ====        and ra, a7, s2
                                                  30'd    9486    : data = 32'h    00279133    ;    //    sll x2 x15 x2      ====        sll sp, a5, sp
                                                  30'd    9487    : data = 32'h    017B24B3    ;    //    slt x9 x22 x23      ====        slt s1, s6, s7
                                                  30'd    9488    : data = 32'h    7D96BE13    ;    //    sltiu x28 x13 2009      ====        sltiu t3, a3, 2009
                                                  30'd    9489    : data = 32'h    016FF633    ;    //    and x12 x31 x22      ====        and a2, t6, s6
                                                  30'd    9490    : data = 32'h    99EC0493    ;    //    addi x9 x24 -1634      ====        addi s1, s8, -1634
                                                  30'd    9491    : data = 32'h    01695313    ;    //    srli x6 x18 22      ====        srli t1, s2, 22
                                                  30'd    9492    : data = 32'h    1529A093    ;    //    slti x1 x19 338      ====        slti ra, s3, 338
                                                  30'd    9493    : data = 32'h    00995EB3    ;    //    srl x29 x18 x9      ====        srl t4, s2, s1
                                                  30'd    9494    : data = 32'h    1ECAF717    ;    //    auipc x14 126127      ====        auipc a4, 126127
                                                  30'd    9495    : data = 32'h    005AD993    ;    //    srli x19 x21 5      ====        srli s3, s5, 5
                                                  30'd    9496    : data = 32'h    0109FFB3    ;    //    and x31 x19 x16      ====        and t6, s3, a6
                                                  30'd    9497    : data = 32'h    DF984813    ;    //    xori x16 x16 -519      ====        xori a6, a6, -519
                                                  30'd    9498    : data = 32'h    01F795B3    ;    //    sll x11 x15 x31      ====        sll a1, a5, t6
                                                  30'd    9499    : data = 32'h    01F35C93    ;    //    srli x25 x6 31      ====        srli s9, t1, 31
                                                  30'd    9500    : data = 32'h    415E5D33    ;    //    sra x26 x28 x21      ====        sra s10, t3, s5
                                                  30'd    9501    : data = 32'h    01FAE3B3    ;    //    or x7 x21 x31      ====        or t2, s5, t6
                                                  30'd    9502    : data = 32'h    AF7EBE37    ;    //    lui x28 718827      ====        lui t3, 718827
                                                  30'd    9503    : data = 32'h    B59AF993    ;    //    andi x19 x21 -1191      ====        andi s3, s5, -1191
                                                  30'd    9504    : data = 32'h    41958C33    ;    //    sub x24 x11 x25      ====        sub s8, a1, s9
                                                  30'd    9505    : data = 32'h    00DA8033    ;    //    add x0 x21 x13      ====        add zero, s5, a3
                                                  30'd    9506    : data = 32'h    01A91DB3    ;    //    sll x27 x18 x26      ====        sll s11, s2, s10
                                                  30'd    9507    : data = 32'h    0032BAB3    ;    //    sltu x21 x5 x3      ====        sltu s5, t0, gp
                                                  30'd    9508    : data = 32'h    8966C593    ;    //    xori x11 x13 -1898      ====        xori a1, a3, -1898
                                                  30'd    9509    : data = 32'h    01B287B3    ;    //    add x15 x5 x27      ====        add a5, t0, s11
                                                  30'd    9510    : data = 32'h    AC822A93    ;    //    slti x21 x4 -1336      ====        slti s5, tp, -1336
                                                  30'd    9511    : data = 32'h    01E45E13    ;    //    srli x28 x8 30      ====        srli t3, s0, 30
                                                  30'd    9512    : data = 32'h    AB5A8B17    ;    //    auipc x22 701864      ====        auipc s6, 701864
                                                  30'd    9513    : data = 32'h    E9F08A13    ;    //    addi x20 x1 -353      ====        addi s4, ra, -353
                                                  30'd    9514    : data = 32'h    4361C137    ;    //    lui x2 275996      ====        lui sp, 275996
                                                  30'd    9515    : data = 32'h    50A74093    ;    //    xori x1 x14 1290      ====        xori ra, a4, 1290
                                                  30'd    9516    : data = 32'h    71910417    ;    //    auipc x8 465168      ====        auipc s0, 465168
                                                  30'd    9517    : data = 32'h    01CB9C13    ;    //    slli x24 x23 28      ====        slli s8, s7, 28
                                                  30'd    9518    : data = 32'h    EF076813    ;    //    ori x16 x14 -272      ====        ori a6, a4, -272
                                                  30'd    9519    : data = 32'h    40A28093    ;    //    addi x1 x5 1034      ====        addi ra, t0, 1034
                                                  30'd    9520    : data = 32'h    0053DE93    ;    //    srli x29 x7 5      ====        srli t4, t2, 5
                                                  30'd    9521    : data = 32'h    24796A93    ;    //    ori x21 x18 583      ====        ori s5, s2, 583
                                                  30'd    9522    : data = 32'h    00A27FB3    ;    //    and x31 x4 x10      ====        and t6, tp, a0
                                                  30'd    9523    : data = 32'h    F7346893    ;    //    ori x17 x8 -141      ====        ori a7, s0, -141
                                                  30'd    9524    : data = 32'h    ECA12793    ;    //    slti x15 x2 -310      ====        slti a5, sp, -310
                                                  30'd    9525    : data = 32'h    00E59633    ;    //    sll x12 x11 x14      ====        sll a2, a1, a4
                                                  30'd    9526    : data = 32'h    01C33DB3    ;    //    sltu x27 x6 x28      ====        sltu s11, t1, t3
                                                  30'd    9527    : data = 32'h    E8CB3B93    ;    //    sltiu x23 x22 -372      ====        sltiu s7, s6, -372
                                                  30'd    9528    : data = 32'h    50BEBD13    ;    //    sltiu x26 x29 1291      ====        sltiu s10, t4, 1291
                                                  30'd    9529    : data = 32'h    00E940B3    ;    //    xor x1 x18 x14      ====        xor ra, s2, a4
                                                  30'd    9530    : data = 32'h    4F230B93    ;    //    addi x23 x6 1266      ====        addi s7, t1, 1266
                                                  30'd    9531    : data = 32'h    F8F75497    ;    //    auipc x9 1019765      ====        auipc s1, 1019765
                                                  30'd    9532    : data = 32'h    4004D013    ;    //    srai x0 x9 0      ====        srai zero, s1, 0
                                                  30'd    9533    : data = 32'h    EB883293    ;    //    sltiu x5 x16 -328      ====        sltiu t0, a6, -328
                                                  30'd    9534    : data = 32'h    CFFE7A93    ;    //    andi x21 x28 -769      ====        andi s5, t3, -769
                                                  30'd    9535    : data = 32'h    008303B3    ;    //    add x7 x6 x8      ====        add t2, t1, s0
                                                  30'd    9536    : data = 32'h    01E6D6B3    ;    //    srl x13 x13 x30      ====        srl a3, a3, t5
                                                  30'd    9537    : data = 32'h    0F0CB493    ;    //    sltiu x9 x25 240      ====        sltiu s1, s9, 240
                                                  30'd    9538    : data = 32'h    40C68633    ;    //    sub x12 x13 x12      ====        sub a2, a3, a2
                                                  30'd    9539    : data = 32'h    83F22997    ;    //    auipc x19 540450      ====        auipc s3, 540450
                                                  30'd    9540    : data = 32'h    00FFB9B3    ;    //    sltu x19 x31 x15      ====        sltu s3, t6, a5
                                                  30'd    9541    : data = 32'h    80000D37    ;    //    lui x26 524288      ====        li s10, 0x80000000 #start riscv_int_numeric_corner_stream_7
                                                  30'd    9542    : data = 32'h    000D0D13    ;    //    addi x26 x26 0      ====        li s10, 0x80000000 #start riscv_int_numeric_corner_stream_7
                                                  30'd    9543    : data = 32'h    800002B7    ;    //    lui x5 524288      ====        li t0, 0x80000000
                                                  30'd    9544    : data = 32'h    00028293    ;    //    addi x5 x5 0      ====        li t0, 0x80000000
                                                  30'd    9545    : data = 32'h    00000593    ;    //    addi x11 x0 0      ====        li a1, 0x0
                                                  30'd    9546    : data = 32'h    800007B7    ;    //    lui x15 524288      ====        li a5, 0x80000000
                                                  30'd    9547    : data = 32'h    00078793    ;    //    addi x15 x15 0      ====        li a5, 0x80000000
                                                  30'd    9548    : data = 32'h    00000893    ;    //    addi x17 x0 0      ====        li a7, 0x0
                                                  30'd    9549    : data = 32'h    1255C337    ;    //    lui x6 75100      ====        li t1, 0x1255b8d1
                                                  30'd    9550    : data = 32'h    8D130313    ;    //    addi x6 x6 -1839      ====        li t1, 0x1255b8d1
                                                  30'd    9551    : data = 32'h    80000DB7    ;    //    lui x27 524288      ====        li s11, 0x80000000
                                                  30'd    9552    : data = 32'h    000D8D93    ;    //    addi x27 x27 0      ====        li s11, 0x80000000
                                                  30'd    9553    : data = 32'h    00000093    ;    //    addi x1 x0 0      ====        li ra, 0x0
                                                  30'd    9554    : data = 32'h    00000A93    ;    //    addi x21 x0 0      ====        li s5, 0x0
                                                  30'd    9555    : data = 32'h    48563637    ;    //    lui x12 296291      ====        li a2, 0x485635b9
                                                  30'd    9556    : data = 32'h    5B960613    ;    //    addi x12 x12 1465      ====        li a2, 0x485635b9
                                                  30'd    9557    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9558    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9559    : data = 32'h    00F88DB3    ;    //    add x27 x17 x15      ====        add s11, a7, a5
                                                  30'd    9560    : data = 32'h    41160333    ;    //    sub x6 x12 x17      ====        sub t1, a2, a7
                                                  30'd    9561    : data = 32'h    00CD87B3    ;    //    add x15 x27 x12      ====        add a5, s11, a2
                                                  30'd    9562    : data = 32'h    14296DB7    ;    //    lui x27 82582      ====        lui s11, 82582
                                                  30'd    9563    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9564    : data = 32'h    35608D13    ;    //    addi x26 x1 854      ====        addi s10, ra, 854
                                                  30'd    9565    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9566    : data = 32'h    D47B5D37    ;    //    lui x26 870325      ====        lui s10, 870325
                                                  30'd    9567    : data = 32'h    D6C30093    ;    //    addi x1 x6 -660      ====        addi ra, t1, -660
                                                  30'd    9568    : data = 32'h    41A88333    ;    //    sub x6 x17 x26      ====        sub t1, a7, s10
                                                  30'd    9569    : data = 32'h    40528D33    ;    //    sub x26 x5 x5      ====        sub s10, t0, t0
                                                  30'd    9570    : data = 32'h    01A60633    ;    //    add x12 x12 x26      ====        add a2, a2, s10
                                                  30'd    9571    : data = 32'h    D5478D13    ;    //    addi x26 x15 -684      ====        addi s10, a5, -684
                                                  30'd    9572    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9573    : data = 32'h    00DC9DB7    ;    //    lui x27 3529      ====        lui s11, 3529
                                                  30'd    9574    : data = 32'h    01AD8AB3    ;    //    add x21 x27 x26      ====        add s5, s11, s10
                                                  30'd    9575    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9576    : data = 32'h    41BD0D33    ;    //    sub x26 x26 x27      ====        sub s10, s10, s11
                                                  30'd    9577    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9578    : data = 32'h    F94C6A97    ;    //    auipc x21 1021126      ====        auipc s5, 1021126
                                                  30'd    9579    : data = 32'h    A2268297    ;    //    auipc x5 664168      ====        auipc t0, 664168
                                                  30'd    9580    : data = 32'h    138020EF    ;    //    jal x1 8504      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_7
                                                  30'd    9581    : data = 32'h    4456E193    ;    //    ori x3 x13 1093      ====        ori gp, a3, 1093
                                                  30'd    9582    : data = 32'h    015086B3    ;    //    add x13 x1 x21      ====        add a3, ra, s5
                                                  30'd    9583    : data = 32'h    01DE1D13    ;    //    slli x26 x28 29      ====        slli s10, t3, 29
                                                  30'd    9584    : data = 32'h    0106D013    ;    //    srli x0 x13 16      ====        srli zero, a3, 16
                                                  30'd    9585    : data = 32'h    40C88133    ;    //    sub x2 x17 x12      ====        sub sp, a7, a2
                                                  30'd    9586    : data = 32'h    C12FE893    ;    //    ori x17 x31 -1006      ====        ori a7, t6, -1006
                                                  30'd    9587    : data = 32'h    0084CC33    ;    //    xor x24 x9 x8      ====        xor s8, s1, s0
                                                  30'd    9588    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9589    : data = 32'h    DC620893    ;    //    addi x17 x4 -570      ====        addi a7, tp, -570
                                                  30'd    9590    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9591    : data = 32'h    49742613    ;    //    slti x12 x8 1175      ====        slti a2, s0, 1175
                                                  30'd    9592    : data = 32'h    0E698113    ;    //    addi x2 x19 230      ====        addi sp, s3, 230
                                                  30'd    9593    : data = 32'h    413082B3    ;    //    sub x5 x1 x19      ====        sub t0, ra, s3
                                                  30'd    9594    : data = 32'h    01EC96B3    ;    //    sll x13 x25 x30      ====        sll a3, s9, t5
                                                  30'd    9595    : data = 32'h    300722B7    ;    //    lui x5 196722      ====        lui t0, 196722
                                                  30'd    9596    : data = 32'h    96CA7C37    ;    //    lui x24 617639      ====        lui s8, 617639
                                                  30'd    9597    : data = 32'h    00269313    ;    //    slli x6 x13 2      ====        slli t1, a3, 2
                                                  30'd    9598    : data = 32'h    01E99D13    ;    //    slli x26 x19 30      ====        slli s10, s3, 30
                                                  30'd    9599    : data = 32'h    01A87833    ;    //    and x16 x16 x26      ====        and a6, a6, s10
                                                  30'd    9600    : data = 32'h    15727913    ;    //    andi x18 x4 343      ====        andi s2, tp, 343
                                                  30'd    9601    : data = 32'h    0122D033    ;    //    srl x0 x5 x18      ====        srl zero, t0, s2
                                                  30'd    9602    : data = 32'h    01BA9693    ;    //    slli x13 x21 27      ====        slli a3, s5, 27
                                                  30'd    9603    : data = 32'h    01BC87B3    ;    //    add x15 x25 x27      ====        add a5, s9, s11
                                                  30'd    9604    : data = 32'h    5C35EC97    ;    //    auipc x25 377694      ====        auipc s9, 377694
                                                  30'd    9605    : data = 32'h    403DD893    ;    //    srai x17 x27 3      ====        srai a7, s11, 3
                                                  30'd    9606    : data = 32'h    6166F713    ;    //    andi x14 x13 1558      ====        andi a4, a3, 1558
                                                  30'd    9607    : data = 32'h    CF0D4613    ;    //    xori x12 x26 -784      ====        xori a2, s10, -784
                                                  30'd    9608    : data = 32'h    419509B3    ;    //    sub x19 x10 x25      ====        sub s3, a0, s9
                                                  30'd    9609    : data = 32'h    010E21B3    ;    //    slt x3 x28 x16      ====        slt gp, t3, a6
                                                  30'd    9610    : data = 32'h    01CBE0B3    ;    //    or x1 x23 x28      ====        or ra, s7, t3
                                                  30'd    9611    : data = 32'h    00FADC13    ;    //    srli x24 x21 15      ====        srli s8, s5, 15
                                                  30'd    9612    : data = 32'h    00796DB3    ;    //    or x27 x18 x7      ====        or s11, s2, t2
                                                  30'd    9613    : data = 32'h    71D32613    ;    //    slti x12 x6 1821      ====        slti a2, t1, 1821
                                                  30'd    9614    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9615    : data = 32'h    00F17733    ;    //    and x14 x2 x15      ====        and a4, sp, a5
                                                  30'd    9616    : data = 32'h    AFF33913    ;    //    sltiu x18 x6 -1281      ====        sltiu s2, t1, -1281
                                                  30'd    9617    : data = 32'h    9F4C2593    ;    //    slti x11 x24 -1548      ====        slti a1, s8, -1548
                                                  30'd    9618    : data = 32'h    0C63E593    ;    //    ori x11 x7 198      ====        ori a1, t2, 198
                                                  30'd    9619    : data = 32'h    B8040B37    ;    //    lui x22 753728      ====        lui s6, 753728
                                                  30'd    9620    : data = 32'h    A5772E13    ;    //    slti x28 x14 -1449      ====        slti t3, a4, -1449
                                                  30'd    9621    : data = 32'h    4085D613    ;    //    srai x12 x11 8      ====        srai a2, a1, 8
                                                  30'd    9622    : data = 32'h    00B45833    ;    //    srl x16 x8 x11      ====        srl a6, s0, a1
                                                  30'd    9623    : data = 32'h    01D4D493    ;    //    srli x9 x9 29      ====        srli s1, s1, 29
                                                  30'd    9624    : data = 32'h    01F49FB3    ;    //    sll x31 x9 x31      ====        sll t6, s1, t6
                                                  30'd    9625    : data = 32'h    013F9113    ;    //    slli x2 x31 19      ====        slli sp, t6, 19
                                                  30'd    9626    : data = 32'h    004DD813    ;    //    srli x16 x27 4      ====        srli a6, s11, 4
                                                  30'd    9627    : data = 32'h    CA566013    ;    //    ori x0 x12 -859      ====        ori zero, a2, -859
                                                  30'd    9628    : data = 32'h    141C8293    ;    //    addi x5 x25 321      ====        addi t0, s9, 321
                                                  30'd    9629    : data = 32'h    001C95B3    ;    //    sll x11 x25 x1      ====        sll a1, s9, ra
                                                  30'd    9630    : data = 32'h    E62CAB93    ;    //    slti x23 x25 -414      ====        slti s7, s9, -414
                                                  30'd    9631    : data = 32'h    01B3DD93    ;    //    srli x27 x7 27      ====        srli s11, t2, 27
                                                  30'd    9632    : data = 32'h    33C48B93    ;    //    addi x23 x9 828      ====        addi s7, s1, 828
                                                  30'd    9633    : data = 32'h    A20E9D37    ;    //    lui x26 663785      ====        lui s10, 663785
                                                  30'd    9634    : data = 32'h    D7B700B7    ;    //    lui x1 883568      ====        lui ra, 883568
                                                  30'd    9635    : data = 32'h    01C15433    ;    //    srl x8 x2 x28      ====        srl s0, sp, t3
                                                  30'd    9636    : data = 32'h    415FD813    ;    //    srai x16 x31 21      ====        srai a6, t6, 21
                                                  30'd    9637    : data = 32'h    67536E13    ;    //    ori x28 x6 1653      ====        ori t3, t1, 1653
                                                  30'd    9638    : data = 32'h    B84C2613    ;    //    slti x12 x24 -1148      ====        slti a2, s8, -1148
                                                  30'd    9639    : data = 32'h    01BE03B3    ;    //    add x7 x28 x27      ====        add t2, t3, s11
                                                  30'd    9640    : data = 32'h    006C6A33    ;    //    or x20 x24 x6      ====        or s4, s8, t1
                                                  30'd    9641    : data = 32'h    01AACA33    ;    //    xor x20 x21 x26      ====        xor s4, s5, s10
                                                  30'd    9642    : data = 32'h    0038BCB3    ;    //    sltu x25 x17 x3      ====        sltu s9, a7, gp
                                                  30'd    9643    : data = 32'h    7B3AB293    ;    //    sltiu x5 x21 1971      ====        sltiu t0, s5, 1971
                                                  30'd    9644    : data = 32'h    00441C33    ;    //    sll x24 x8 x4      ====        sll s8, s0, tp
                                                  30'd    9645    : data = 32'h    01607433    ;    //    and x8 x0 x22      ====        and s0, zero, s6
                                                  30'd    9646    : data = 32'h    01F25693    ;    //    srli x13 x4 31      ====        srli a3, tp, 31
                                                  30'd    9647    : data = 32'h    7A824D13    ;    //    xori x26 x4 1960      ====        xori s10, tp, 1960
                                                  30'd    9648    : data = 32'h    01FD83B3    ;    //    add x7 x27 x31      ====        add t2, s11, t6
                                                  30'd    9649    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9650    : data = 32'h    41E4DD13    ;    //    srai x26 x9 30      ====        srai s10, s1, 30
                                                  30'd    9651    : data = 32'h    3ED3EE13    ;    //    ori x28 x7 1005      ====        ori t3, t2, 1005
                                                  30'd    9652    : data = 32'h    00A424B3    ;    //    slt x9 x8 x10      ====        slt s1, s0, a0
                                                  30'd    9653    : data = 32'h    CC4EBE93    ;    //    sltiu x29 x29 -828      ====        sltiu t4, t4, -828
                                                  30'd    9654    : data = 32'h    00D05E93    ;    //    srli x29 x0 13      ====        srli t4, zero, 13
                                                  30'd    9655    : data = 32'h    78A2F013    ;    //    andi x0 x5 1930      ====        andi zero, t0, 1930
                                                  30'd    9656    : data = 32'h    003B07B3    ;    //    add x15 x22 x3      ====        add a5, s6, gp
                                                  30'd    9657    : data = 32'h    4AF1E693    ;    //    ori x13 x3 1199      ====        ori a3, gp, 1199
                                                  30'd    9658    : data = 32'h    01DD8CB3    ;    //    add x25 x27 x29      ====        add s9, s11, t4
                                                  30'd    9659    : data = 32'h    00D73B33    ;    //    sltu x22 x14 x13      ====        sltu s6, a4, a3
                                                  30'd    9660    : data = 32'h    01C3D6B3    ;    //    srl x13 x7 x28      ====        srl a3, t2, t3
                                                  30'd    9661    : data = 32'h    0036BB33    ;    //    sltu x22 x13 x3      ====        sltu s6, a3, gp
                                                  30'd    9662    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9663    : data = 32'h    DDE9DD37    ;    //    lui x26 908957      ====        lui s10, 908957
                                                  30'd    9664    : data = 32'h    DDEC7013    ;    //    andi x0 x24 -546      ====        andi zero, s8, -546
                                                  30'd    9665    : data = 32'h    403356B3    ;    //    sra x13 x6 x3      ====        sra a3, t1, gp
                                                  30'd    9666    : data = 32'h    A9A209B7    ;    //    lui x19 694816      ====        lui s3, 694816
                                                  30'd    9667    : data = 32'h    01F0FA33    ;    //    and x20 x1 x31      ====        and s4, ra, t6
                                                  30'd    9668    : data = 32'h    00BE9FB3    ;    //    sll x31 x29 x11      ====        sll t6, t4, a1
                                                  30'd    9669    : data = 32'h    0065DC93    ;    //    srli x25 x11 6      ====        srli s9, a1, 6
                                                  30'd    9670    : data = 32'h    01AC9493    ;    //    slli x9 x25 26      ====        slli s1, s9, 26
                                                  30'd    9671    : data = 32'h    4097DE93    ;    //    srai x29 x15 9      ====        srai t4, a5, 9
                                                  30'd    9672    : data = 32'h    00151EB3    ;    //    sll x29 x10 x1      ====        sll t4, a0, ra
                                                  30'd    9673    : data = 32'h    0081DD33    ;    //    srl x26 x3 x8      ====        srl s10, gp, s0
                                                  30'd    9674    : data = 32'h    B20EC993    ;    //    xori x19 x29 -1248      ====        xori s3, t4, -1248
                                                  30'd    9675    : data = 32'h    417C0DB3    ;    //    sub x27 x24 x23      ====        sub s11, s8, s7
                                                  30'd    9676    : data = 32'h    9C36F993    ;    //    andi x19 x13 -1597      ====        andi s3, a3, -1597
                                                  30'd    9677    : data = 32'h    01EC1033    ;    //    sll x0 x24 x30      ====        sll zero, s8, t5
                                                  30'd    9678    : data = 32'h    0148F4B3    ;    //    and x9 x17 x20      ====        and s1, a7, s4
                                                  30'd    9679    : data = 32'h    B30C7593    ;    //    andi x11 x24 -1232      ====        andi a1, s8, -1232
                                                  30'd    9680    : data = 32'h    F4FFE593    ;    //    ori x11 x31 -177      ====        ori a1, t6, -177
                                                  30'd    9681    : data = 32'h    015A42B3    ;    //    xor x5 x20 x21      ====        xor t0, s4, s5
                                                  30'd    9682    : data = 32'h    4123DA13    ;    //    srai x20 x7 18      ====        srai s4, t2, 18
                                                  30'd    9683    : data = 32'h    40015B33    ;    //    sra x22 x2 x0      ====        sra s6, sp, zero
                                                  30'd    9684    : data = 32'h    01589A33    ;    //    sll x20 x17 x21      ====        sll s4, a7, s5
                                                  30'd    9685    : data = 32'h    01B02433    ;    //    slt x8 x0 x27      ====        slt s0, zero, s11
                                                  30'd    9686    : data = 32'h    01A364B3    ;    //    or x9 x6 x26      ====        or s1, t1, s10
                                                  30'd    9687    : data = 32'h    0005ECB3    ;    //    or x25 x11 x0      ====        or s9, a1, zero
                                                  30'd    9688    : data = 32'h    00B03433    ;    //    sltu x8 x0 x11      ====        sltu s0, zero, a1
                                                  30'd    9689    : data = 32'h    0B35C297    ;    //    auipc x5 45916      ====        auipc t0, 45916
                                                  30'd    9690    : data = 32'h    017B4D33    ;    //    xor x26 x22 x23      ====        xor s10, s6, s7
                                                  30'd    9691    : data = 32'h    00314EB3    ;    //    xor x29 x2 x3      ====        xor t4, sp, gp
                                                  30'd    9692    : data = 32'h    012C9A93    ;    //    slli x21 x25 18      ====        slli s5, s9, 18
                                                  30'd    9693    : data = 32'h    88D8AC93    ;    //    slti x25 x17 -1907      ====        slti s9, a7, -1907
                                                  30'd    9694    : data = 32'h    0027FE33    ;    //    and x28 x15 x2      ====        and t3, a5, sp
                                                  30'd    9695    : data = 32'h    01F73433    ;    //    sltu x8 x14 x31      ====        sltu s0, a4, t6
                                                  30'd    9696    : data = 32'h    BEF56897    ;    //    auipc x17 782166      ====        auipc a7, 782166
                                                  30'd    9697    : data = 32'h    B01EE093    ;    //    ori x1 x29 -1279      ====        ori ra, t4, -1279
                                                  30'd    9698    : data = 32'h    015F9E33    ;    //    sll x28 x31 x21      ====        sll t3, t6, s5
                                                  30'd    9699    : data = 32'h    000EF833    ;    //    and x16 x29 x0      ====        and a6, t4, zero
                                                  30'd    9700    : data = 32'h    0094E1B3    ;    //    or x3 x9 x9      ====        or gp, s1, s1
                                                  30'd    9701    : data = 32'h    001A45B3    ;    //    xor x11 x20 x1      ====        xor a1, s4, ra
                                                  30'd    9702    : data = 32'h    40B85293    ;    //    srai x5 x16 11      ====        srai t0, a6, 11
                                                  30'd    9703    : data = 32'h    14DC2817    ;    //    auipc x16 85442      ====        auipc a6, 85442
                                                  30'd    9704    : data = 32'h    00CEE7B3    ;    //    or x15 x29 x12      ====        or a5, t4, a2
                                                  30'd    9705    : data = 32'h    00C01BB3    ;    //    sll x23 x0 x12      ====        sll s7, zero, a2
                                                  30'd    9706    : data = 32'h    00D507B3    ;    //    add x15 x10 x13      ====        add a5, a0, a3
                                                  30'd    9707    : data = 32'h    01275AB3    ;    //    srl x21 x14 x18      ====        srl s5, a4, s2
                                                  30'd    9708    : data = 32'h    0117F4B3    ;    //    and x9 x15 x17      ====        and s1, a5, a7
                                                  30'd    9709    : data = 32'h    407D0833    ;    //    sub x16 x26 x7      ====        sub a6, s10, t2
                                                  30'd    9710    : data = 32'h    00122633    ;    //    slt x12 x4 x1      ====        slt a2, tp, ra
                                                  30'd    9711    : data = 32'h    40CC8CB3    ;    //    sub x25 x25 x12      ====        sub s9, s9, a2
                                                  30'd    9712    : data = 32'h    01E975B3    ;    //    and x11 x18 x30      ====        and a1, s2, t5
                                                  30'd    9713    : data = 32'h    1E58BB93    ;    //    sltiu x23 x17 485      ====        sltiu s7, a7, 485
                                                  30'd    9714    : data = 32'h    A732DE37    ;    //    lui x28 684845      ====        lui t3, 684845
                                                  30'd    9715    : data = 32'h    01F5DBB3    ;    //    srl x23 x11 x31      ====        srl s7, a1, t6
                                                  30'd    9716    : data = 32'h    3E7E5A37    ;    //    lui x20 255973      ====        lui s4, 255973
                                                  30'd    9717    : data = 32'h    548D3D13    ;    //    sltiu x26 x26 1352      ====        sltiu s10, s10, 1352
                                                  30'd    9718    : data = 32'h    01B19093    ;    //    slli x1 x3 27      ====        slli ra, gp, 27
                                                  30'd    9719    : data = 32'h    010E1393    ;    //    slli x7 x28 16      ====        slli t2, t3, 16
                                                  30'd    9720    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9721    : data = 32'h    013D3DB3    ;    //    sltu x27 x26 x19      ====        sltu s11, s10, s3
                                                  30'd    9722    : data = 32'h    00A5C433    ;    //    xor x8 x11 x10      ====        xor s0, a1, a0
                                                  30'd    9723    : data = 32'h    8B5CB013    ;    //    sltiu x0 x25 -1867      ====        sltiu zero, s9, -1867
                                                  30'd    9724    : data = 32'h    01A05593    ;    //    srli x11 x0 26      ====        srli a1, zero, 26
                                                  30'd    9725    : data = 32'h    41775493    ;    //    srai x9 x14 23      ====        srai s1, a4, 23
                                                  30'd    9726    : data = 32'h    013B1993    ;    //    slli x19 x22 19      ====        slli s3, s6, 19
                                                  30'd    9727    : data = 32'h    3238A393    ;    //    slti x7 x17 803      ====        slti t2, a7, 803
                                                  30'd    9728    : data = 32'h    42ED4B13    ;    //    xori x22 x26 1070      ====        xori s6, s10, 1070
                                                  30'd    9729    : data = 32'h    EDB09337    ;    //    lui x6 973577      ====        lui t1, 973577
                                                  30'd    9730    : data = 32'h    ECA2AF93    ;    //    slti x31 x5 -310      ====        slti t6, t0, -310
                                                  30'd    9731    : data = 32'h    00DF9433    ;    //    sll x8 x31 x13      ====        sll s0, t6, a3
                                                  30'd    9732    : data = 32'h    019F4EB3    ;    //    xor x29 x30 x25      ====        xor t4, t5, s9
                                                  30'd    9733    : data = 32'h    01549733    ;    //    sll x14 x9 x21      ====        sll a4, s1, s5
                                                  30'd    9734    : data = 32'h    EAFC2B37    ;    //    lui x22 962498      ====        lui s6, 962498
                                                  30'd    9735    : data = 32'h    E1798293    ;    //    addi x5 x19 -489      ====        addi t0, s3, -489
                                                  30'd    9736    : data = 32'h    1417C1B7    ;    //    lui x3 82300      ====        lui gp, 82300
                                                  30'd    9737    : data = 32'h    015FB833    ;    //    sltu x16 x31 x21      ====        sltu a6, t6, s5
                                                  30'd    9738    : data = 32'h    36CF3713    ;    //    sltiu x14 x30 876      ====        sltiu a4, t5, 876
                                                  30'd    9739    : data = 32'h    00968B33    ;    //    add x22 x13 x9      ====        add s6, a3, s1
                                                  30'd    9740    : data = 32'h    01165C13    ;    //    srli x24 x12 17      ====        srli s8, a2, 17
                                                  30'd    9741    : data = 32'h    FBFA8113    ;    //    addi x2 x21 -65      ====        addi sp, s5, -65
                                                  30'd    9742    : data = 32'h    01ED0EB3    ;    //    add x29 x26 x30      ====        add t4, s10, t5
                                                  30'd    9743    : data = 32'h    412B0E33    ;    //    sub x28 x22 x18      ====        sub t3, s6, s2
                                                  30'd    9744    : data = 32'h    4C580E13    ;    //    addi x28 x16 1221      ====        addi t3, a6, 1221
                                                  30'd    9745    : data = 32'h    016F7C93    ;    //    andi x25 x30 22      ====        andi s9, t5, 22
                                                  30'd    9746    : data = 32'h    00970033    ;    //    add x0 x14 x9      ====        add zero, a4, s1
                                                  30'd    9747    : data = 32'h    0136F133    ;    //    and x2 x13 x19      ====        and sp, a3, s3
                                                  30'd    9748    : data = 32'h    0178CFB3    ;    //    xor x31 x17 x23      ====        xor t6, a7, s7
                                                  30'd    9749    : data = 32'h    0184B133    ;    //    sltu x2 x9 x24      ====        sltu sp, s1, s8
                                                  30'd    9750    : data = 32'h    F42DAB93    ;    //    slti x23 x27 -190      ====        slti s7, s11, -190
                                                  30'd    9751    : data = 32'h    9452A613    ;    //    slti x12 x5 -1723      ====        slti a2, t0, -1723
                                                  30'd    9752    : data = 32'h    41C98E33    ;    //    sub x28 x19 x28      ====        sub t3, s3, t3
                                                  30'd    9753    : data = 32'h    4137D713    ;    //    srai x14 x15 19      ====        srai a4, a5, 19
                                                  30'd    9754    : data = 32'h    00A0C133    ;    //    xor x2 x1 x10      ====        xor sp, ra, a0
                                                  30'd    9755    : data = 32'h    F6274913    ;    //    xori x18 x14 -158      ====        xori s2, a4, -158
                                                  30'd    9756    : data = 32'h    00C249B3    ;    //    xor x19 x4 x12      ====        xor s3, tp, a2
                                                  30'd    9757    : data = 32'h    01235833    ;    //    srl x16 x6 x18      ====        srl a6, t1, s2
                                                  30'd    9758    : data = 32'h    4136DCB3    ;    //    sra x25 x13 x19      ====        sra s9, a3, s3
                                                  30'd    9759    : data = 32'h    005EEFB3    ;    //    or x31 x29 x5      ====        or t6, t4, t0
                                                  30'd    9760    : data = 32'h    00B27A33    ;    //    and x20 x4 x11      ====        and s4, tp, a1
                                                  30'd    9761    : data = 32'h    45E7D737    ;    //    lui x14 286333      ====        lui a4, 286333
                                                  30'd    9762    : data = 32'h    4117D0B3    ;    //    sra x1 x15 x17      ====        sra ra, a5, a7
                                                  30'd    9763    : data = 32'h    00475413    ;    //    srli x8 x14 4      ====        srli s0, a4, 4
                                                  30'd    9764    : data = 32'h    412E8A33    ;    //    sub x20 x29 x18      ====        sub s4, t4, s2
                                                  30'd    9765    : data = 32'h    D976E593    ;    //    ori x11 x13 -617      ====        ori a1, a3, -617
                                                  30'd    9766    : data = 32'h    0026F9B3    ;    //    and x19 x13 x2      ====        and s3, a3, sp
                                                  30'd    9767    : data = 32'h    01ADD193    ;    //    srli x3 x27 26      ====        srli gp, s11, 26
                                                  30'd    9768    : data = 32'h    00348733    ;    //    add x14 x9 x3      ====        add a4, s1, gp
                                                  30'd    9769    : data = 32'h    1B47B693    ;    //    sltiu x13 x15 436      ====        sltiu a3, a5, 436
                                                  30'd    9770    : data = 32'h    7A744813    ;    //    xori x16 x8 1959      ====        xori a6, s0, 1959
                                                  30'd    9771    : data = 32'h    41097E17    ;    //    auipc x28 266391      ====        auipc t3, 266391
                                                  30'd    9772    : data = 32'h    410B5393    ;    //    srai x7 x22 16      ====        srai t2, s6, 16
                                                  30'd    9773    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9774    : data = 32'h    01A15693    ;    //    srli x13 x2 26      ====        srli a3, sp, 26
                                                  30'd    9775    : data = 32'h    51B89A37    ;    //    lui x20 334729      ====        lui s4, 334729
                                                  30'd    9776    : data = 32'h    37798C93    ;    //    addi x25 x19 887      ====        addi s9, s3, 887
                                                  30'd    9777    : data = 32'h    019B5C13    ;    //    srli x24 x22 25      ====        srli s8, s6, 25
                                                  30'd    9778    : data = 32'h    0060DB93    ;    //    srli x23 x1 6      ====        srli s7, ra, 6
                                                  30'd    9779    : data = 32'h    00A3F033    ;    //    and x0 x7 x10      ====        and zero, t2, a0
                                                  30'd    9780    : data = 32'h    055B0A37    ;    //    lui x20 21936      ====        lui s4, 21936
                                                  30'd    9781    : data = 32'h    001670B3    ;    //    and x1 x12 x1      ====        and ra, a2, ra
                                                  30'd    9782    : data = 32'h    F0258613    ;    //    addi x12 x11 -254      ====        addi a2, a1, -254
                                                  30'd    9783    : data = 32'h    011191B3    ;    //    sll x3 x3 x17      ====        sll gp, gp, a7
                                                  30'd    9784    : data = 32'h    01DADA13    ;    //    srli x20 x21 29      ====        srli s4, s5, 29
                                                  30'd    9785    : data = 32'h    0175DD13    ;    //    srli x26 x11 23      ====        srli s10, a1, 23
                                                  30'd    9786    : data = 32'h    9378BE17    ;    //    auipc x28 604043      ====        auipc t3, 604043
                                                  30'd    9787    : data = 32'h    9F644C13    ;    //    xori x24 x8 -1546      ====        xori s8, s0, -1546
                                                  30'd    9788    : data = 32'h    40BEDA33    ;    //    sra x20 x29 x11      ====        sra s4, t4, a1
                                                  30'd    9789    : data = 32'h    4330CB17    ;    //    auipc x22 275212      ====        auipc s6, 275212
                                                  30'd    9790    : data = 32'h    4181DEB3    ;    //    sra x29 x3 x24      ====        sra t4, gp, s8
                                                  30'd    9791    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9792    : data = 32'h    001763B3    ;    //    or x7 x14 x1      ====        or t2, a4, ra
                                                  30'd    9793    : data = 32'h    01C8A1B3    ;    //    slt x3 x17 x28      ====        slt gp, a7, t3
                                                  30'd    9794    : data = 32'h    412AD7B3    ;    //    sra x15 x21 x18      ====        sra a5, s5, s2
                                                  30'd    9795    : data = 32'h    0061D033    ;    //    srl x0 x3 x6      ====        srl zero, gp, t1
                                                  30'd    9796    : data = 32'h    0106B833    ;    //    sltu x16 x13 x16      ====        sltu a6, a3, a6
                                                  30'd    9797    : data = 32'h    01D5C033    ;    //    xor x0 x11 x29      ====        xor zero, a1, t4
                                                  30'd    9798    : data = 32'h    402E5013    ;    //    srai x0 x28 2      ====        srai zero, t3, 2
                                                  30'd    9799    : data = 32'h    0008B6B3    ;    //    sltu x13 x17 x0      ====        sltu a3, a7, zero
                                                  30'd    9800    : data = 32'h    40950BB3    ;    //    sub x23 x10 x9      ====        sub s7, a0, s1
                                                  30'd    9801    : data = 32'h    0153C4B3    ;    //    xor x9 x7 x21      ====        xor s1, t2, s5
                                                  30'd    9802    : data = 32'h    64047B13    ;    //    andi x22 x8 1600      ====        andi s6, s0, 1600
                                                  30'd    9803    : data = 32'h    00F5A033    ;    //    slt x0 x11 x15      ====        slt zero, a1, a5
                                                  30'd    9804    : data = 32'h    416F04B3    ;    //    sub x9 x30 x22      ====        sub s1, t5, s6
                                                  30'd    9805    : data = 32'h    13070C93    ;    //    addi x25 x14 304      ====        addi s9, a4, 304
                                                  30'd    9806    : data = 32'h    01B79393    ;    //    slli x7 x15 27      ====        slli t2, a5, 27
                                                  30'd    9807    : data = 32'h    F8DE7593    ;    //    andi x11 x28 -115      ====        andi a1, t3, -115
                                                  30'd    9808    : data = 32'h    FBD42713    ;    //    slti x14 x8 -67      ====        slti a4, s0, -67
                                                  30'd    9809    : data = 32'h    4043DA93    ;    //    srai x21 x7 4      ====        srai s5, t2, 4
                                                  30'd    9810    : data = 32'h    5B8DAE13    ;    //    slti x28 x27 1464      ====        slti t3, s11, 1464
                                                  30'd    9811    : data = 32'h    00F796B3    ;    //    sll x13 x15 x15      ====        sll a3, a5, a5
                                                  30'd    9812    : data = 32'h    40D40E33    ;    //    sub x28 x8 x13      ====        sub t3, s0, a3
                                                  30'd    9813    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9814    : data = 32'h    ADC63893    ;    //    sltiu x17 x12 -1316      ====        sltiu a7, a2, -1316
                                                  30'd    9815    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9816    : data = 32'h    86220E13    ;    //    addi x28 x4 -1950      ====        addi t3, tp, -1950
                                                  30'd    9817    : data = 32'h    00A9FD33    ;    //    and x26 x19 x10      ====        and s10, s3, a0
                                                  30'd    9818    : data = 32'h    0191CEB3    ;    //    xor x29 x3 x25      ====        xor t4, gp, s9
                                                  30'd    9819    : data = 32'h    3C036D93    ;    //    ori x27 x6 960      ====        ori s11, t1, 960
                                                  30'd    9820    : data = 32'h    002ED713    ;    //    srli x14 x29 2      ====        srli a4, t4, 2
                                                  30'd    9821    : data = 32'h    00DAA933    ;    //    slt x18 x21 x13      ====        slt s2, s5, a3
                                                  30'd    9822    : data = 32'h    011A0FB3    ;    //    add x31 x20 x17      ====        add t6, s4, a7
                                                  30'd    9823    : data = 32'h    01E35433    ;    //    srl x8 x6 x30      ====        srl s0, t1, t5
                                                  30'd    9824    : data = 32'h    00034E13    ;    //    xori x28 x6 0      ====        xori t3, t1, 0
                                                  30'd    9825    : data = 32'h    01DE4C33    ;    //    xor x24 x28 x29      ====        xor s8, t3, t4
                                                  30'd    9826    : data = 32'h    DFADEB13    ;    //    ori x22 x27 -518      ====        ori s6, s11, -518
                                                  30'd    9827    : data = 32'h    11754713    ;    //    xori x14 x10 279      ====        xori a4, a0, 279
                                                  30'd    9828    : data = 32'h    75E4EA13    ;    //    ori x20 x9 1886      ====        ori s4, s1, 1886
                                                  30'd    9829    : data = 32'h    2647CE13    ;    //    xori x28 x15 612      ====        xori t3, a5, 612
                                                  30'd    9830    : data = 32'h    B1243193    ;    //    sltiu x3 x8 -1262      ====        sltiu gp, s0, -1262
                                                  30'd    9831    : data = 32'h    01D95933    ;    //    srl x18 x18 x29      ====        srl s2, s2, t4
                                                  30'd    9832    : data = 32'h    01F94B33    ;    //    xor x22 x18 x31      ====        xor s6, s2, t6
                                                  30'd    9833    : data = 32'h    008117B3    ;    //    sll x15 x2 x8      ====        sll a5, sp, s0
                                                  30'd    9834    : data = 32'h    475D7B13    ;    //    andi x22 x26 1141      ====        andi s6, s10, 1141
                                                  30'd    9835    : data = 32'h    014996B3    ;    //    sll x13 x19 x20      ====        sll a3, s3, s4
                                                  30'd    9836    : data = 32'h    1397A693    ;    //    slti x13 x15 313      ====        slti a3, a5, 313
                                                  30'd    9837    : data = 32'h    1A50EA13    ;    //    ori x20 x1 421      ====        ori s4, ra, 421
                                                  30'd    9838    : data = 32'h    05FF8D93    ;    //    addi x27 x31 95      ====        addi s11, t6, 95
                                                  30'd    9839    : data = 32'h    D926AE17    ;    //    auipc x28 889450      ====        auipc t3, 889450
                                                  30'd    9840    : data = 32'h    79EF3937    ;    //    lui x18 499443      ====        lui s2, 499443
                                                  30'd    9841    : data = 32'h    FEE9F397    ;    //    auipc x7 1044127      ====        auipc t2, 1044127
                                                  30'd    9842    : data = 32'h    000D1833    ;    //    sll x16 x26 x0      ====        sll a6, s10, zero
                                                  30'd    9843    : data = 32'h    018908B3    ;    //    add x17 x18 x24      ====        add a7, s2, s8
                                                  30'd    9844    : data = 32'h    1A643F97    ;    //    auipc x31 108099      ====        auipc t6, 108099
                                                  30'd    9845    : data = 32'h    01F77633    ;    //    and x12 x14 x31      ====        and a2, a4, t6
                                                  30'd    9846    : data = 32'h    0331A313    ;    //    slti x6 x3 51      ====        slti t1, gp, 51
                                                  30'd    9847    : data = 32'h    010B15B3    ;    //    sll x11 x22 x16      ====        sll a1, s6, a6
                                                  30'd    9848    : data = 32'h    01F2D733    ;    //    srl x14 x5 x31      ====        srl a4, t0, t6
                                                  30'd    9849    : data = 32'h    4158DB13    ;    //    srai x22 x17 21      ====        srai s6, a7, 21
                                                  30'd    9850    : data = 32'h    502FA797    ;    //    auipc x15 328442      ====        auipc a5, 328442
                                                  30'd    9851    : data = 32'h    41A4DBB3    ;    //    sra x23 x9 x26      ====        sra s7, s1, s10
                                                  30'd    9852    : data = 32'h    DA9B7B93    ;    //    andi x23 x22 -599      ====        andi s7, s6, -599
                                                  30'd    9853    : data = 32'h    417C5B33    ;    //    sra x22 x24 x23      ====        sra s6, s8, s7
                                                  30'd    9854    : data = 32'h    41D03A13    ;    //    sltiu x20 x0 1053      ====        sltiu s4, zero, 1053
                                                  30'd    9855    : data = 32'h    01A59E13    ;    //    slli x28 x11 26      ====        slli t3, a1, 26
                                                  30'd    9856    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9857    : data = 32'h    977A2E17    ;    //    auipc x28 620450      ====        auipc t3, 620450
                                                  30'd    9858    : data = 32'h    01E4B033    ;    //    sltu x0 x9 x30      ====        sltu zero, s1, t5
                                                  30'd    9859    : data = 32'h    414A86B3    ;    //    sub x13 x21 x20      ====        sub a3, s5, s4
                                                  30'd    9860    : data = 32'h    41DC8433    ;    //    sub x8 x25 x29      ====        sub s0, s9, t4
                                                  30'd    9861    : data = 32'h    00447D33    ;    //    and x26 x8 x4      ====        and s10, s0, tp
                                                  30'd    9862    : data = 32'h    01E13833    ;    //    sltu x16 x2 x30      ====        sltu a6, sp, t5
                                                  30'd    9863    : data = 32'h    41E10D33    ;    //    sub x26 x2 x30      ====        sub s10, sp, t5
                                                  30'd    9864    : data = 32'h    01229F93    ;    //    slli x31 x5 18      ====        slli t6, t0, 18
                                                  30'd    9865    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9866    : data = 32'h    A986C113    ;    //    xori x2 x13 -1384      ====        xori sp, a3, -1384
                                                  30'd    9867    : data = 32'h    01F5C333    ;    //    xor x6 x11 x31      ====        xor t1, a1, t6
                                                  30'd    9868    : data = 32'h    0013B733    ;    //    sltu x14 x7 x1      ====        sltu a4, t2, ra
                                                  30'd    9869    : data = 32'h    0172CBB3    ;    //    xor x23 x5 x23      ====        xor s7, t0, s7
                                                  30'd    9870    : data = 32'h    67712593    ;    //    slti x11 x2 1655      ====        slti a1, sp, 1655
                                                  30'd    9871    : data = 32'h    A8297297    ;    //    auipc x5 688791      ====        auipc t0, 688791
                                                  30'd    9872    : data = 32'h    8AA58D93    ;    //    addi x27 x11 -1878      ====        addi s11, a1, -1878
                                                  30'd    9873    : data = 32'h    40A05CB3    ;    //    sra x25 x0 x10      ====        sra s9, zero, a0
                                                  30'd    9874    : data = 32'h    01FB0A33    ;    //    add x20 x22 x31      ====        add s4, s6, t6
                                                  30'd    9875    : data = 32'h    5AF832B7    ;    //    lui x5 372611      ====        lui t0, 372611
                                                  30'd    9876    : data = 32'h    303CB097    ;    //    auipc x1 197579      ====        auipc ra, 197579
                                                  30'd    9877    : data = 32'h    A9A87A93    ;    //    andi x21 x16 -1382      ====        andi s5, a6, -1382
                                                  30'd    9878    : data = 32'h    00E0BB33    ;    //    sltu x22 x1 x14      ====        sltu s6, ra, a4
                                                  30'd    9879    : data = 32'h    01F5E733    ;    //    or x14 x11 x31      ====        or a4, a1, t6
                                                  30'd    9880    : data = 32'h    000412B3    ;    //    sll x5 x8 x0      ====        sll t0, s0, zero
                                                  30'd    9881    : data = 32'h    414F83B3    ;    //    sub x7 x31 x20      ====        sub t2, t6, s4
                                                  30'd    9882    : data = 32'h    00141C33    ;    //    sll x24 x8 x1      ====        sll s8, s0, ra
                                                  30'd    9883    : data = 32'h    005CACB3    ;    //    slt x25 x25 x5      ====        slt s9, s9, t0
                                                  30'd    9884    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9885    : data = 32'h    215C4393    ;    //    xori x7 x24 533      ====        xori t2, s8, 533
                                                  30'd    9886    : data = 32'h    B0374997    ;    //    auipc x19 721780      ====        auipc s3, 721780
                                                  30'd    9887    : data = 32'h    0169D013    ;    //    srli x0 x19 22      ====        srli zero, s3, 22
                                                  30'd    9888    : data = 32'h    408D56B3    ;    //    sra x13 x26 x8      ====        sra a3, s10, s0
                                                  30'd    9889    : data = 32'h    829F2713    ;    //    slti x14 x30 -2007      ====        slti a4, t5, -2007
                                                  30'd    9890    : data = 32'h    00CDBD33    ;    //    sltu x26 x27 x12      ====        sltu s10, s11, a2
                                                  30'd    9891    : data = 32'h    725BF313    ;    //    andi x6 x23 1829      ====        andi t1, s7, 1829
                                                  30'd    9892    : data = 32'h    41C45A13    ;    //    srai x20 x8 28      ====        srai s4, s0, 28
                                                  30'd    9893    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9894    : data = 32'h    417ADE33    ;    //    sra x28 x21 x23      ====        sra t3, s5, s7
                                                  30'd    9895    : data = 32'h    41CDD413    ;    //    srai x8 x27 28      ====        srai s0, s11, 28
                                                  30'd    9896    : data = 32'h    01455BB3    ;    //    srl x23 x10 x20      ====        srl s7, a0, s4
                                                  30'd    9897    : data = 32'h    011D1C13    ;    //    slli x24 x26 17      ====        slli s8, s10, 17
                                                  30'd    9898    : data = 32'h    0139F1B3    ;    //    and x3 x19 x19      ====        and gp, s3, s3
                                                  30'd    9899    : data = 32'h    41ED5033    ;    //    sra x0 x26 x30      ====        sra zero, s10, t5
                                                  30'd    9900    : data = 32'h    C5DDF593    ;    //    andi x11 x27 -931      ====        andi a1, s11, -931
                                                  30'd    9901    : data = 32'h    006A9833    ;    //    sll x16 x21 x6      ====        sll a6, s5, t1
                                                  30'd    9902    : data = 32'h    D020E913    ;    //    ori x18 x1 -766      ====        ori s2, ra, -766
                                                  30'd    9903    : data = 32'h    018FCAB3    ;    //    xor x21 x31 x24      ====        xor s5, t6, s8
                                                  30'd    9904    : data = 32'h    4054D033    ;    //    sra x0 x9 x5      ====        sra zero, s1, t0
                                                  30'd    9905    : data = 32'h    01E5ED33    ;    //    or x26 x11 x30      ====        or s10, a1, t5
                                                  30'd    9906    : data = 32'h    00539493    ;    //    slli x9 x7 5      ====        slli s1, t2, 5
                                                  30'd    9907    : data = 32'h    003BA4B3    ;    //    slt x9 x23 x3      ====        slt s1, s7, gp
                                                  30'd    9908    : data = 32'h    910CE093    ;    //    ori x1 x25 -1776      ====        ori ra, s9, -1776
                                                  30'd    9909    : data = 32'h    01D3C933    ;    //    xor x18 x7 x29      ====        xor s2, t2, t4
                                                  30'd    9910    : data = 32'h    0009BDB3    ;    //    sltu x27 x19 x0      ====        sltu s11, s3, zero
                                                  30'd    9911    : data = 32'h    015F65B3    ;    //    or x11 x30 x21      ====        or a1, t5, s5
                                                  30'd    9912    : data = 32'h    0190EFB3    ;    //    or x31 x1 x25      ====        or t6, ra, s9
                                                  30'd    9913    : data = 32'h    014E1033    ;    //    sll x0 x28 x20      ====        sll zero, t3, s4
                                                  30'd    9914    : data = 32'h    407E8DB3    ;    //    sub x27 x29 x7      ====        sub s11, t4, t2
                                                  30'd    9915    : data = 32'h    00AB35B3    ;    //    sltu x11 x22 x10      ====        sltu a1, s6, a0
                                                  30'd    9916    : data = 32'h    00EC9CB3    ;    //    sll x25 x25 x14      ====        sll s9, s9, a4
                                                  30'd    9917    : data = 32'h    00C9D7B3    ;    //    srl x15 x19 x12      ====        srl a5, s3, a2
                                                  30'd    9918    : data = 32'h    015D5633    ;    //    srl x12 x26 x21      ====        srl a2, s10, s5
                                                  30'd    9919    : data = 32'h    228CAF93    ;    //    slti x31 x25 552      ====        slti t6, s9, 552
                                                  30'd    9920    : data = 32'h    01CFE8B3    ;    //    or x17 x31 x28      ====        or a7, t6, t3
                                                  30'd    9921    : data = 32'h    415F8433    ;    //    sub x8 x31 x21      ====        sub s0, t6, s5
                                                  30'd    9922    : data = 32'h    41875F93    ;    //    srai x31 x14 24      ====        srai t6, a4, 24
                                                  30'd    9923    : data = 32'h    0085DAB3    ;    //    srl x21 x11 x8      ====        srl s5, a1, s0
                                                  30'd    9924    : data = 32'h    DB297613    ;    //    andi x12 x18 -590      ====        andi a2, s2, -590
                                                  30'd    9925    : data = 32'h    1687AAB7    ;    //    lui x21 92282      ====        lui s5, 92282
                                                  30'd    9926    : data = 32'h    0179B433    ;    //    sltu x8 x19 x23      ====        sltu s0, s3, s7
                                                  30'd    9927    : data = 32'h    0120DD13    ;    //    srli x26 x1 18      ====        srli s10, ra, 18
                                                  30'd    9928    : data = 32'h    23BDBD13    ;    //    sltiu x26 x27 571      ====        sltiu s10, s11, 571
                                                  30'd    9929    : data = 32'h    012C0033    ;    //    add x0 x24 x18      ====        add zero, s8, s2
                                                  30'd    9930    : data = 32'h    014216B3    ;    //    sll x13 x4 x20      ====        sll a3, tp, s4
                                                  30'd    9931    : data = 32'h    00205BB3    ;    //    srl x23 x0 x2      ====        srl s7, zero, sp
                                                  30'd    9932    : data = 32'h    D5457F93    ;    //    andi x31 x10 -684      ====        andi t6, a0, -684
                                                  30'd    9933    : data = 32'h    726BCA93    ;    //    xori x21 x23 1830      ====        xori s5, s7, 1830
                                                  30'd    9934    : data = 32'h    5651AE13    ;    //    slti x28 x3 1381      ====        slti t3, gp, 1381
                                                  30'd    9935    : data = 32'h    AC094613    ;    //    xori x12 x18 -1344      ====        xori a2, s2, -1344
                                                  30'd    9936    : data = 32'h    019A14B3    ;    //    sll x9 x20 x25      ====        sll s1, s4, s9
                                                  30'd    9937    : data = 32'h    005CACB3    ;    //    slt x25 x25 x5      ====        slt s9, s9, t0
                                                  30'd    9938    : data = 32'h    007A5113    ;    //    srli x2 x20 7      ====        srli sp, s4, 7
                                                  30'd    9939    : data = 32'h    D173AA13    ;    //    slti x20 x7 -745      ====        slti s4, t2, -745
                                                  30'd    9940    : data = 32'h    0177F5B3    ;    //    and x11 x15 x23      ====        and a1, a5, s7
                                                  30'd    9941    : data = 32'h    00C4D793    ;    //    srli x15 x9 12      ====        srli a5, s1, 12
                                                  30'd    9942    : data = 32'h    00D925B3    ;    //    slt x11 x18 x13      ====        slt a1, s2, a3
                                                  30'd    9943    : data = 32'h    4093DD93    ;    //    srai x27 x7 9      ====        srai s11, t2, 9
                                                  30'd    9944    : data = 32'h    40D55093    ;    //    srai x1 x10 13      ====        srai ra, a0, 13
                                                  30'd    9945    : data = 32'h    01445793    ;    //    srli x15 x8 20      ====        srli a5, s0, 20
                                                  30'd    9946    : data = 32'h    00DC96B3    ;    //    sll x13 x25 x13      ====        sll a3, s9, a3
                                                  30'd    9947    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9948    : data = 32'h    010955B3    ;    //    srl x11 x18 x16      ====        srl a1, s2, a6
                                                  30'd    9949    : data = 32'h    48A39D17    ;    //    auipc x26 297529      ====        auipc s10, 297529
                                                  30'd    9950    : data = 32'h    EB2CEC93    ;    //    ori x25 x25 -334      ====        ori s9, s9, -334
                                                  30'd    9951    : data = 32'h    00A8CDB3    ;    //    xor x27 x17 x10      ====        xor s11, a7, a0
                                                  30'd    9952    : data = 32'h    015C5EB3    ;    //    srl x29 x24 x21      ====        srl t4, s8, s5
                                                  30'd    9953    : data = 32'h    1CFF6193    ;    //    ori x3 x30 463      ====        ori gp, t5, 463
                                                  30'd    9954    : data = 32'h    C8ECA413    ;    //    slti x8 x25 -882      ====        slti s0, s9, -882
                                                  30'd    9955    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9956    : data = 32'h    01DD6DB3    ;    //    or x27 x26 x29      ====        or s11, s10, t4
                                                  30'd    9957    : data = 32'h    0165D633    ;    //    srl x12 x11 x22      ====        srl a2, a1, s6
                                                  30'd    9958    : data = 32'h    014E86B3    ;    //    add x13 x29 x20      ====        add a3, t4, s4
                                                  30'd    9959    : data = 32'h    C93D3893    ;    //    sltiu x17 x26 -877      ====        sltiu a7, s10, -877
                                                  30'd    9960    : data = 32'h    01D70E33    ;    //    add x28 x14 x29      ====        add t3, a4, t4
                                                  30'd    9961    : data = 32'h    20600D17    ;    //    auipc x26 132608      ====        auipc s10, 132608
                                                  30'd    9962    : data = 32'h    4C35BE93    ;    //    sltiu x29 x11 1219      ====        sltiu t4, a1, 1219
                                                  30'd    9963    : data = 32'h    4810B093    ;    //    sltiu x1 x1 1153      ====        sltiu ra, ra, 1153
                                                  30'd    9964    : data = 32'h    7C5CB713    ;    //    sltiu x14 x25 1989      ====        sltiu a4, s9, 1989
                                                  30'd    9965    : data = 32'h    DA9A8B93    ;    //    addi x23 x21 -599      ====        addi s7, s5, -599
                                                  30'd    9966    : data = 32'h    405FDA93    ;    //    srai x21 x31 5      ====        srai s5, t6, 5
                                                  30'd    9967    : data = 32'h    01F05EB3    ;    //    srl x29 x0 x31      ====        srl t4, zero, t6
                                                  30'd    9968    : data = 32'h    015BEC33    ;    //    or x24 x23 x21      ====        or s8, s7, s5
                                                  30'd    9969    : data = 32'h    41A85013    ;    //    srai x0 x16 26      ====        srai zero, a6, 26
                                                  30'd    9970    : data = 32'h    00C87A33    ;    //    and x20 x16 x12      ====        and s4, a6, a2
                                                  30'd    9971    : data = 32'h    589EA993    ;    //    slti x19 x29 1417      ====        slti s3, t4, 1417
                                                  30'd    9972    : data = 32'h    40C9D393    ;    //    srai x7 x19 12      ====        srai t2, s3, 12
                                                  30'd    9973    : data = 32'h    41A45CB3    ;    //    sra x25 x8 x26      ====        sra s9, s0, s10
                                                  30'd    9974    : data = 32'h    0059B733    ;    //    sltu x14 x19 x5      ====        sltu a4, s3, t0
                                                  30'd    9975    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    9976    : data = 32'h    D93F8BB7    ;    //    lui x23 889848      ====        lui s7, 889848
                                                  30'd    9977    : data = 32'h    6C803613    ;    //    sltiu x12 x0 1736      ====        sltiu a2, zero, 1736
                                                  30'd    9978    : data = 32'h    A5A39397    ;    //    auipc x7 678457      ====        auipc t2, 678457
                                                  30'd    9979    : data = 32'h    FF9DC313    ;    //    xori x6 x27 -7      ====        xori t1, s11, -7
                                                  30'd    9980    : data = 32'h    8B4925B7    ;    //    lui x11 570514      ====        lui a1, 570514
                                                  30'd    9981    : data = 32'h    DC60C5B7    ;    //    lui x11 902668      ====        lui a1, 902668
                                                  30'd    9982    : data = 32'h    DBED2B37    ;    //    lui x22 900818      ====        lui s6, 900818
                                                  30'd    9983    : data = 32'h    A54BDA37    ;    //    lui x20 677053      ====        lui s4, 677053
                                                  30'd    9984    : data = 32'h    00FE12B3    ;    //    sll x5 x28 x15      ====        sll t0, t3, a5
                                                  30'd    9985    : data = 32'h    01A4DA13    ;    //    srli x20 x9 26      ====        srli s4, s1, 26
                                                  30'd    9986    : data = 32'h    167AC313    ;    //    xori x6 x21 359      ====        xori t1, s5, 359
                                                  30'd    9987    : data = 32'h    19BE0D13    ;    //    addi x26 x28 411      ====        addi s10, t3, 411
                                                  30'd    9988    : data = 32'h    37C8F793    ;    //    andi x15 x17 892      ====        andi a5, a7, 892
                                                  30'd    9989    : data = 32'h    0173EDB3    ;    //    or x27 x7 x23      ====        or s11, t2, s7
                                                  30'd    9990    : data = 32'h    40245913    ;    //    srai x18 x8 2      ====        srai s2, s0, 2
                                                  30'd    9991    : data = 32'h    0186EEB3    ;    //    or x29 x13 x24      ====        or t4, a3, s8
                                                  30'd    9992    : data = 32'h    001BB933    ;    //    sltu x18 x23 x1      ====        sltu s2, s7, ra
                                                  30'd    9993    : data = 32'h    4154DE13    ;    //    srai x28 x9 21      ====        srai t3, s1, 21
                                                  30'd    9994    : data = 32'h    AF057B13    ;    //    andi x22 x10 -1296      ====        andi s6, a0, -1296
                                                  30'd    9995    : data = 32'h    B4E04B13    ;    //    xori x22 x0 -1202      ====        xori s6, zero, -1202
                                                  30'd    9996    : data = 32'h    000C5833    ;    //    srl x16 x24 x0      ====        srl a6, s8, zero
                                                  30'd    9997    : data = 32'h    41175B13    ;    //    srai x22 x14 17      ====        srai s6, a4, 17
                                                  30'd    9998    : data = 32'h    004C7AB3    ;    //    and x21 x24 x4      ====        and s5, s8, tp
                                                  30'd    9999    : data = 32'h    0057BA33    ;    //    sltu x20 x15 x5      ====        sltu s4, a5, t0
                                                  30'd    10000    : data = 32'h    01343D33    ;    //    sltu x26 x8 x19      ====        sltu s10, s0, s3
                                                  30'd    10001    : data = 32'h    6EE4B813    ;    //    sltiu x16 x9 1774      ====        sltiu a6, s1, 1774
                                                  30'd    10002    : data = 32'h    41B7DB33    ;    //    sra x22 x15 x27      ====        sra s6, a5, s11
                                                  30'd    10003    : data = 32'h    01FC5CB3    ;    //    srl x25 x24 x31      ====        srl s9, s8, t6
                                                  30'd    10004    : data = 32'h    001ADEB3    ;    //    srl x29 x21 x1      ====        srl t4, s5, ra
                                                  30'd    10005    : data = 32'h    4D5ED5B7    ;    //    lui x11 316909      ====        lui a1, 316909
                                                  30'd    10006    : data = 32'h    416D86B3    ;    //    sub x13 x27 x22      ====        sub a3, s11, s6
                                                  30'd    10007    : data = 32'h    40135093    ;    //    srai x1 x6 1      ====        srai ra, t1, 1
                                                  30'd    10008    : data = 32'h    017E90B3    ;    //    sll x1 x29 x23      ====        sll ra, t4, s7
                                                  30'd    10009    : data = 32'h    40A7D593    ;    //    srai x11 x15 10      ====        srai a1, a5, 10
                                                  30'd    10010    : data = 32'h    18BCF593    ;    //    andi x11 x25 395      ====        andi a1, s9, 395
                                                  30'd    10011    : data = 32'h    00B79013    ;    //    slli x0 x15 11      ====        slli zero, a5, 11
                                                  30'd    10012    : data = 32'h    000BDE93    ;    //    srli x29 x23 0      ====        srli t4, s7, 0
                                                  30'd    10013    : data = 32'h    415456B3    ;    //    sra x13 x8 x21      ====        sra a3, s0, s5
                                                  30'd    10014    : data = 32'h    01EB6333    ;    //    or x6 x22 x30      ====        or t1, s6, t5
                                                  30'd    10015    : data = 32'h    41B35E33    ;    //    sra x28 x6 x27      ====        sra t3, t1, s11
                                                  30'd    10016    : data = 32'h    40BB8B33    ;    //    sub x22 x23 x11      ====        sub s6, s7, a1
                                                  30'd    10017    : data = 32'h    550CF693    ;    //    andi x13 x25 1360      ====        andi a3, s9, 1360
                                                  30'd    10018    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10019    : data = 32'h    00541713    ;    //    slli x14 x8 5      ====        slli a4, s0, 5
                                                  30'd    10020    : data = 32'h    00C15E13    ;    //    srli x28 x2 12      ====        srli t3, sp, 12
                                                  30'd    10021    : data = 32'h    00B11593    ;    //    slli x11 x2 11      ====        slli a1, sp, 11
                                                  30'd    10022    : data = 32'h    01736C33    ;    //    or x24 x6 x23      ====        or s8, t1, s7
                                                  30'd    10023    : data = 32'h    EA3E8113    ;    //    addi x2 x29 -349      ====        addi sp, t4, -349
                                                  30'd    10024    : data = 32'h    408C8A33    ;    //    sub x20 x25 x8      ====        sub s4, s9, s0
                                                  30'd    10025    : data = 32'h    00584833    ;    //    xor x16 x16 x5      ====        xor a6, a6, t0
                                                  30'd    10026    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10027    : data = 32'h    C6729DB7    ;    //    lui x27 812841      ====        lui s11, 812841
                                                  30'd    10028    : data = 32'h    1AB3EB13    ;    //    ori x22 x7 427      ====        ori s6, t2, 427
                                                  30'd    10029    : data = 32'h    00755133    ;    //    srl x2 x10 x7      ====        srl sp, a0, t2
                                                  30'd    10030    : data = 32'h    01FF3733    ;    //    sltu x14 x30 x31      ====        sltu a4, t5, t6
                                                  30'd    10031    : data = 32'h    01F881B3    ;    //    add x3 x17 x31      ====        add gp, a7, t6
                                                  30'd    10032    : data = 32'h    41D0D913    ;    //    srai x18 x1 29      ====        srai s2, ra, 29
                                                  30'd    10033    : data = 32'h    006BB5B3    ;    //    sltu x11 x23 x6      ====        sltu a1, s7, t1
                                                  30'd    10034    : data = 32'h    40EC8733    ;    //    sub x14 x25 x14      ====        sub a4, s9, a4
                                                  30'd    10035    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10036    : data = 32'h    01D582B3    ;    //    add x5 x11 x29      ====        add t0, a1, t4
                                                  30'd    10037    : data = 32'h    00846EB3    ;    //    or x29 x8 x8      ====        or t4, s0, s0
                                                  30'd    10038    : data = 32'h    1586B613    ;    //    sltiu x12 x13 344      ====        sltiu a2, a3, 344
                                                  30'd    10039    : data = 32'h    00CF7DB3    ;    //    and x27 x30 x12      ====        and s11, t5, a2
                                                  30'd    10040    : data = 32'h    408A5C33    ;    //    sra x24 x20 x8      ====        sra s8, s4, s0
                                                  30'd    10041    : data = 32'h    3E583A93    ;    //    sltiu x21 x16 997      ====        sltiu s5, a6, 997
                                                  30'd    10042    : data = 32'h    00511C33    ;    //    sll x24 x2 x5      ====        sll s8, sp, t0
                                                  30'd    10043    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10044    : data = 32'h    D534EAB7    ;    //    lui x21 873294      ====        lui s5, 873294
                                                  30'd    10045    : data = 32'h    004D8133    ;    //    add x2 x27 x4      ====        add sp, s11, tp
                                                  30'd    10046    : data = 32'h    00DDD893    ;    //    srli x17 x27 13      ====        srli a7, s11, 13
                                                  30'd    10047    : data = 32'h    B8B50B13    ;    //    addi x22 x10 -1141      ====        addi s6, a0, -1141
                                                  30'd    10048    : data = 32'h    4160DAB3    ;    //    sra x21 x1 x22      ====        sra s5, ra, s6
                                                  30'd    10049    : data = 32'h    86E8CB13    ;    //    xori x22 x17 -1938      ====        xori s6, a7, -1938
                                                  30'd    10050    : data = 32'h    0018AE33    ;    //    slt x28 x17 x1      ====        slt t3, a7, ra
                                                  30'd    10051    : data = 32'h    8CACA613    ;    //    slti x12 x25 -1846      ====        slti a2, s9, -1846
                                                  30'd    10052    : data = 32'h    90E9BCB7    ;    //    lui x25 593563      ====        lui s9, 593563
                                                  30'd    10053    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10054    : data = 32'h    00545E93    ;    //    srli x29 x8 5      ====        srli t4, s0, 5
                                                  30'd    10055    : data = 32'h    40C4D5B3    ;    //    sra x11 x9 x12      ====        sra a1, s1, a2
                                                  30'd    10056    : data = 32'h    01CDE7B3    ;    //    or x15 x27 x28      ====        or a5, s11, t3
                                                  30'd    10057    : data = 32'h    008AA833    ;    //    slt x16 x21 x8      ====        slt a6, s5, s0
                                                  30'd    10058    : data = 32'h    01AE1793    ;    //    slli x15 x28 26      ====        slli a5, t3, 26
                                                  30'd    10059    : data = 32'h    2C923E93    ;    //    sltiu x29 x4 713      ====        sltiu t4, tp, 713
                                                  30'd    10060    : data = 32'h    019C5113    ;    //    srli x2 x24 25      ====        srli sp, s8, 25
                                                  30'd    10061    : data = 32'h    41FD5713    ;    //    srai x14 x26 31      ====        srai a4, s10, 31
                                                  30'd    10062    : data = 32'h    A543B1B7    ;    //    lui x3 676923      ====        lui gp, 676923
                                                  30'd    10063    : data = 32'h    01B7D713    ;    //    srli x14 x15 27      ====        srli a4, a5, 27
                                                  30'd    10064    : data = 32'h    65936393    ;    //    ori x7 x6 1625      ====        ori t2, t1, 1625
                                                  30'd    10065    : data = 32'h    01B08833    ;    //    add x16 x1 x27      ====        add a6, ra, s11
                                                  30'd    10066    : data = 32'h    6771DA97    ;    //    auipc x21 423709      ====        auipc s5, 423709
                                                  30'd    10067    : data = 32'h    5E0B7693    ;    //    andi x13 x22 1504      ====        andi a3, s6, 1504
                                                  30'd    10068    : data = 32'h    46716D13    ;    //    ori x26 x2 1127      ====        ori s10, sp, 1127
                                                  30'd    10069    : data = 32'h    0F756A13    ;    //    ori x20 x10 247      ====        ori s4, a0, 247
                                                  30'd    10070    : data = 32'h    19E1B593    ;    //    sltiu x11 x3 414      ====        sltiu a1, gp, 414
                                                  30'd    10071    : data = 32'h    2339B593    ;    //    sltiu x11 x19 563      ====        sltiu a1, s3, 563
                                                  30'd    10072    : data = 32'h    007B9613    ;    //    slli x12 x23 7      ====        slli a2, s7, 7
                                                  30'd    10073    : data = 32'h    413FD393    ;    //    srai x7 x31 19      ====        srai t2, t6, 19
                                                  30'd    10074    : data = 32'h    23F51A37    ;    //    lui x20 147281      ====        lui s4, 147281
                                                  30'd    10075    : data = 32'h    0102E033    ;    //    or x0 x5 x16      ====        or zero, t0, a6
                                                  30'd    10076    : data = 32'h    001FE3B3    ;    //    or x7 x31 x1      ====        or t2, t6, ra
                                                  30'd    10077    : data = 32'h    00921D93    ;    //    slli x27 x4 9      ====        slli s11, tp, 9
                                                  30'd    10078    : data = 32'h    00F7B933    ;    //    sltu x18 x15 x15      ====        sltu s2, a5, a5
                                                  30'd    10079    : data = 32'h    65014B93    ;    //    xori x23 x2 1616      ====        xori s7, sp, 1616
                                                  30'd    10080    : data = 32'h    A9293613    ;    //    sltiu x12 x18 -1390      ====        sltiu a2, s2, -1390
                                                  30'd    10081    : data = 32'h    4014D333    ;    //    sra x6 x9 x1      ====        sra t1, s1, ra
                                                  30'd    10082    : data = 32'h    01452EB3    ;    //    slt x29 x10 x20      ====        slt t4, a0, s4
                                                  30'd    10083    : data = 32'h    005BC8B3    ;    //    xor x17 x23 x5      ====        xor a7, s7, t0
                                                  30'd    10084    : data = 32'h    011DD433    ;    //    srl x8 x27 x17      ====        srl s0, s11, a7
                                                  30'd    10085    : data = 32'h    401FD3B3    ;    //    sra x7 x31 x1      ====        sra t2, t6, ra
                                                  30'd    10086    : data = 32'h    01F451B3    ;    //    srl x3 x8 x31      ====        srl gp, s0, t6
                                                  30'd    10087    : data = 32'h    41B15E33    ;    //    sra x28 x2 x27      ====        sra t3, sp, s11
                                                  30'd    10088    : data = 32'h    20549A17    ;    //    auipc x20 132425      ====        auipc s4, 132425
                                                  30'd    10089    : data = 32'h    7F570713    ;    //    addi x14 x14 2037      ====        addi a4, a4, 2037
                                                  30'd    10090    : data = 32'h    01911313    ;    //    slli x6 x2 25      ====        slli t1, sp, 25
                                                  30'd    10091    : data = 32'h    00EFD6B3    ;    //    srl x13 x31 x14      ====        srl a3, t6, a4
                                                  30'd    10092    : data = 32'h    2200F693    ;    //    andi x13 x1 544      ====        andi a3, ra, 544
                                                  30'd    10093    : data = 32'h    CE253B37    ;    //    lui x22 844371      ====        lui s6, 844371
                                                  30'd    10094    : data = 32'h    003F1DB3    ;    //    sll x27 x30 x3      ====        sll s11, t5, gp
                                                  30'd    10095    : data = 32'h    326D7293    ;    //    andi x5 x26 806      ====        andi t0, s10, 806
                                                  30'd    10096    : data = 32'h    E753F437    ;    //    lui x8 947519      ====        lui s0, 947519
                                                  30'd    10097    : data = 32'h    DC8A4413    ;    //    xori x8 x20 -568      ====        xori s0, s4, -568
                                                  30'd    10098    : data = 32'h    01626133    ;    //    or x2 x4 x22      ====        or sp, tp, s6
                                                  30'd    10099    : data = 32'h    01D93EB3    ;    //    sltu x29 x18 x29      ====        sltu t4, s2, t4
                                                  30'd    10100    : data = 32'h    4038D693    ;    //    srai x13 x17 3      ====        srai a3, a7, 3
                                                  30'd    10101    : data = 32'h    004C8E33    ;    //    add x28 x25 x4      ====        add t3, s9, tp
                                                  30'd    10102    : data = 32'h    A0608E13    ;    //    addi x28 x1 -1530      ====        addi t3, ra, -1530
                                                  30'd    10103    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10104    : data = 32'h    002DC0B3    ;    //    xor x1 x27 x2      ====        xor ra, s11, sp
                                                  30'd    10105    : data = 32'h    C1D58193    ;    //    addi x3 x11 -995      ====        addi gp, a1, -995
                                                  30'd    10106    : data = 32'h    007B1693    ;    //    slli x13 x22 7      ====        slli a3, s6, 7
                                                  30'd    10107    : data = 32'h    406ED113    ;    //    srai x2 x29 6      ====        srai sp, t4, 6
                                                  30'd    10108    : data = 32'h    41835FB3    ;    //    sra x31 x6 x24      ====        sra t6, t1, s8
                                                  30'd    10109    : data = 32'h    00BAD5B3    ;    //    srl x11 x21 x11      ====        srl a1, s5, a1
                                                  30'd    10110    : data = 32'h    005B9893    ;    //    slli x17 x23 5      ====        slli a7, s7, 5
                                                  30'd    10111    : data = 32'h    1F30AE13    ;    //    slti x28 x1 499      ====        slti t3, ra, 499
                                                  30'd    10112    : data = 32'h    01E19833    ;    //    sll x16 x3 x30      ====        sll a6, gp, t5
                                                  30'd    10113    : data = 32'h    D06D46B7    ;    //    lui x13 853716      ====        lui a3, 853716
                                                  30'd    10114    : data = 32'h    1B036A13    ;    //    ori x20 x6 432      ====        ori s4, t1, 432
                                                  30'd    10115    : data = 32'h    0064AA33    ;    //    slt x20 x9 x6      ====        slt s4, s1, t1
                                                  30'd    10116    : data = 32'h    01D9DA33    ;    //    srl x20 x19 x29      ====        srl s4, s3, t4
                                                  30'd    10117    : data = 32'h    00E14AB3    ;    //    xor x21 x2 x14      ====        xor s5, sp, a4
                                                  30'd    10118    : data = 32'h    418FDB33    ;    //    sra x22 x31 x24      ====        sra s6, t6, s8
                                                  30'd    10119    : data = 32'h    01221913    ;    //    slli x18 x4 18      ====        slli s2, tp, 18
                                                  30'd    10120    : data = 32'h    0A48C393    ;    //    xori x7 x17 164      ====        xori t2, a7, 164
                                                  30'd    10121    : data = 32'h    0096D5B3    ;    //    srl x11 x13 x9      ====        srl a1, a3, s1
                                                  30'd    10122    : data = 32'h    008E2EB3    ;    //    slt x29 x28 x8      ====        slt t4, t3, s0
                                                  30'd    10123    : data = 32'h    01ED7733    ;    //    and x14 x26 x30      ====        and a4, s10, t5
                                                  30'd    10124    : data = 32'h    409A0033    ;    //    sub x0 x20 x9      ====        sub zero, s4, s1
                                                  30'd    10125    : data = 32'h    413F5F93    ;    //    srai x31 x30 19      ====        srai t6, t5, 19
                                                  30'd    10126    : data = 32'h    70AC6A93    ;    //    ori x21 x24 1802      ====        ori s5, s8, 1802
                                                  30'd    10127    : data = 32'h    0162BFB3    ;    //    sltu x31 x5 x22      ====        sltu t6, t0, s6
                                                  30'd    10128    : data = 32'h    C9B0C717    ;    //    auipc x14 826124      ====        auipc a4, 826124
                                                  30'd    10129    : data = 32'h    007774B3    ;    //    and x9 x14 x7      ====        and s1, a4, t2
                                                  30'd    10130    : data = 32'h    FBE68293    ;    //    addi x5 x13 -66      ====        addi t0, a3, -66
                                                  30'd    10131    : data = 32'h    001F5713    ;    //    srli x14 x30 1      ====        srli a4, t5, 1
                                                  30'd    10132    : data = 32'h    87A9AF93    ;    //    slti x31 x19 -1926      ====        slti t6, s3, -1926
                                                  30'd    10133    : data = 32'h    00BDD693    ;    //    srli x13 x27 11      ====        srli a3, s11, 11
                                                  30'd    10134    : data = 32'h    EF29D417    ;    //    auipc x8 979613      ====        auipc s0, 979613
                                                  30'd    10135    : data = 32'h    7BA69297    ;    //    auipc x5 506473      ====        auipc t0, 506473
                                                  30'd    10136    : data = 32'h    40BD56B3    ;    //    sra x13 x26 x11      ====        sra a3, s10, a1
                                                  30'd    10137    : data = 32'h    40F15C13    ;    //    srai x24 x2 15      ====        srai s8, sp, 15
                                                  30'd    10138    : data = 32'h    E5E1C893    ;    //    xori x17 x3 -418      ====        xori a7, gp, -418
                                                  30'd    10139    : data = 32'h    0148A6B3    ;    //    slt x13 x17 x20      ====        slt a3, a7, s4
                                                  30'd    10140    : data = 32'h    01806593    ;    //    ori x11 x0 24      ====        ori a1, zero, 24
                                                  30'd    10141    : data = 32'h    00CC1AB3    ;    //    sll x21 x24 x12      ====        sll s5, s8, a2
                                                  30'd    10142    : data = 32'h    40B25433    ;    //    sra x8 x4 x11      ====        sra s0, tp, a1
                                                  30'd    10143    : data = 32'h    63F6E917    ;    //    auipc x18 409454      ====        auipc s2, 409454
                                                  30'd    10144    : data = 32'h    001A1913    ;    //    slli x18 x20 1      ====        slli s2, s4, 1
                                                  30'd    10145    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10146    : data = 32'h    0199A0B3    ;    //    slt x1 x19 x25      ====        slt ra, s3, s9
                                                  30'd    10147    : data = 32'h    007C5293    ;    //    srli x5 x24 7      ====        srli t0, s8, 7
                                                  30'd    10148    : data = 32'h    4134D6B3    ;    //    sra x13 x9 x19      ====        sra a3, s1, s3
                                                  30'd    10149    : data = 32'h    00A2FCB3    ;    //    and x25 x5 x10      ====        and s9, t0, a0
                                                  30'd    10150    : data = 32'h    173C7A93    ;    //    andi x21 x24 371      ====        andi s5, s8, 371
                                                  30'd    10151    : data = 32'h    0120FFB3    ;    //    and x31 x1 x18      ====        and t6, ra, s2
                                                  30'd    10152    : data = 32'h    D12CE013    ;    //    ori x0 x25 -750      ====        ori zero, s9, -750
                                                  30'd    10153    : data = 32'h    00298EB3    ;    //    add x29 x19 x2      ====        add t4, s3, sp
                                                  30'd    10154    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10155    : data = 32'h    012450B3    ;    //    srl x1 x8 x18      ====        srl ra, s0, s2
                                                  30'd    10156    : data = 32'h    90F97293    ;    //    andi x5 x18 -1777      ====        andi t0, s2, -1777
                                                  30'd    10157    : data = 32'h    01561C13    ;    //    slli x24 x12 21      ====        slli s8, a2, 21
                                                  30'd    10158    : data = 32'h    1284D897    ;    //    auipc x17 75853      ====        auipc a7, 75853
                                                  30'd    10159    : data = 32'h    011F9593    ;    //    slli x11 x31 17      ====        slli a1, t6, 17
                                                  30'd    10160    : data = 32'h    41BCDC13    ;    //    srai x24 x25 27      ====        srai s8, s9, 27
                                                  30'd    10161    : data = 32'h    007BAC33    ;    //    slt x24 x23 x7      ====        slt s8, s7, t2
                                                  30'd    10162    : data = 32'h    018B1393    ;    //    slli x7 x22 24      ====        slli t2, s6, 24
                                                  30'd    10163    : data = 32'h    006F9A93    ;    //    slli x21 x31 6      ====        slli s5, t6, 6
                                                  30'd    10164    : data = 32'h    6A835B37    ;    //    lui x22 436277      ====        lui s6, 436277
                                                  30'd    10165    : data = 32'h    4178DD93    ;    //    srai x27 x17 23      ====        srai s11, a7, 23
                                                  30'd    10166    : data = 32'h    009CB933    ;    //    sltu x18 x25 x9      ====        sltu s2, s9, s1
                                                  30'd    10167    : data = 32'h    7871E413    ;    //    ori x8 x3 1927      ====        ori s0, gp, 1927
                                                  30'd    10168    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10169    : data = 32'h    41F38313    ;    //    addi x6 x7 1055      ====        addi t1, t2, 1055
                                                  30'd    10170    : data = 32'h    5BC37313    ;    //    andi x6 x6 1468      ====        andi t1, t1, 1468
                                                  30'd    10171    : data = 32'h    8AFE8893    ;    //    addi x17 x29 -1873      ====        addi a7, t4, -1873
                                                  30'd    10172    : data = 32'h    D83F3613    ;    //    sltiu x12 x30 -637      ====        sltiu a2, t5, -637
                                                  30'd    10173    : data = 32'h    01D93CB3    ;    //    sltu x25 x18 x29      ====        sltu s9, s2, t4
                                                  30'd    10174    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10175    : data = 32'h    40115433    ;    //    sra x8 x2 x1      ====        sra s0, sp, ra
                                                  30'd    10176    : data = 32'h    33AF2293    ;    //    slti x5 x30 826      ====        slti t0, t5, 826
                                                  30'd    10177    : data = 32'h    41E85593    ;    //    srai x11 x16 30      ====        srai a1, a6, 30
                                                  30'd    10178    : data = 32'h    006E6CB3    ;    //    or x25 x28 x6      ====        or s9, t3, t1
                                                  30'd    10179    : data = 32'h    001E1293    ;    //    slli x5 x28 1      ====        slli t0, t3, 1
                                                  30'd    10180    : data = 32'h    F212A713    ;    //    slti x14 x5 -223      ====        slti a4, t0, -223
                                                  30'd    10181    : data = 32'h    01685313    ;    //    srli x6 x16 22      ====        srli t1, a6, 22
                                                  30'd    10182    : data = 32'h    DF8FA113    ;    //    slti x2 x31 -520      ====        slti sp, t6, -520
                                                  30'd    10183    : data = 32'h    F4121717    ;    //    auipc x14 999713      ====        auipc a4, 999713
                                                  30'd    10184    : data = 32'h    005E0733    ;    //    add x14 x28 x5      ====        add a4, t3, t0
                                                  30'd    10185    : data = 32'h    00EEFAB3    ;    //    and x21 x29 x14      ====        and s5, t4, a4
                                                  30'd    10186    : data = 32'h    00B03733    ;    //    sltu x14 x0 x11      ====        sltu a4, zero, a1
                                                  30'd    10187    : data = 32'h    00F0FDB3    ;    //    and x27 x1 x15      ====        and s11, ra, a5
                                                  30'd    10188    : data = 32'h    16578D93    ;    //    addi x27 x15 357      ====        addi s11, a5, 357
                                                  30'd    10189    : data = 32'h    00FA07B3    ;    //    add x15 x20 x15      ====        add a5, s4, a5
                                                  30'd    10190    : data = 32'h    01A4C133    ;    //    xor x2 x9 x26      ====        xor sp, s1, s10
                                                  30'd    10191    : data = 32'h    01C24CB3    ;    //    xor x25 x4 x28      ====        xor s9, tp, t3
                                                  30'd    10192    : data = 32'h    95E08E13    ;    //    addi x28 x1 -1698      ====        addi t3, ra, -1698
                                                  30'd    10193    : data = 32'h    CCD2BC13    ;    //    sltiu x24 x5 -819      ====        sltiu s8, t0, -819
                                                  30'd    10194    : data = 32'h    41475AB3    ;    //    sra x21 x14 x20      ====        sra s5, a4, s4
                                                  30'd    10195    : data = 32'h    01FD1433    ;    //    sll x8 x26 x31      ====        sll s0, s10, t6
                                                  30'd    10196    : data = 32'h    00C388B3    ;    //    add x17 x7 x12      ====        add a7, t2, a2
                                                  30'd    10197    : data = 32'h    00630033    ;    //    add x0 x6 x6      ====        add zero, t1, t1
                                                  30'd    10198    : data = 32'h    896F7B93    ;    //    andi x23 x30 -1898      ====        andi s7, t5, -1898
                                                  30'd    10199    : data = 32'h    01529FB3    ;    //    sll x31 x5 x21      ====        sll t6, t0, s5
                                                  30'd    10200    : data = 32'h    00325713    ;    //    srli x14 x4 3      ====        srli a4, tp, 3
                                                  30'd    10201    : data = 32'h    01BA1713    ;    //    slli x14 x20 27      ====        slli a4, s4, 27
                                                  30'd    10202    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10203    : data = 32'h    40CB04B3    ;    //    sub x9 x22 x12      ====        sub s1, s6, a2
                                                  30'd    10204    : data = 32'h    93BEBA13    ;    //    sltiu x20 x29 -1733      ====        sltiu s4, t4, -1733
                                                  30'd    10205    : data = 32'h    CDFA2013    ;    //    slti x0 x20 -801      ====        slti zero, s4, -801
                                                  30'd    10206    : data = 32'h    4122D6B3    ;    //    sra x13 x5 x18      ====        sra a3, t0, s2
                                                  30'd    10207    : data = 32'h    AB75BD13    ;    //    sltiu x26 x11 -1353      ====        sltiu s10, a1, -1353
                                                  30'd    10208    : data = 32'h    409D5EB3    ;    //    sra x29 x26 x9      ====        sra t4, s10, s1
                                                  30'd    10209    : data = 32'h    300C1717    ;    //    auipc x14 196801      ====        auipc a4, 196801
                                                  30'd    10210    : data = 32'h    0067A033    ;    //    slt x0 x15 x6      ====        slt zero, a5, t1
                                                  30'd    10211    : data = 32'h    410A5793    ;    //    srai x15 x20 16      ====        srai a5, s4, 16
                                                  30'd    10212    : data = 32'h    01E02B33    ;    //    slt x22 x0 x30      ====        slt s6, zero, t5
                                                  30'd    10213    : data = 32'h    016A8E33    ;    //    add x28 x21 x22      ====        add t3, s5, s6
                                                  30'd    10214    : data = 32'h    77296D93    ;    //    ori x27 x18 1906      ====        ori s11, s2, 1906
                                                  30'd    10215    : data = 32'h    405E5793    ;    //    srai x15 x28 5      ====        srai a5, t3, 5
                                                  30'd    10216    : data = 32'h    011877B3    ;    //    and x15 x16 x17      ====        and a5, a6, a7
                                                  30'd    10217    : data = 32'h    01F0CB33    ;    //    xor x22 x1 x31      ====        xor s6, ra, t6
                                                  30'd    10218    : data = 32'h    8BA0AD93    ;    //    slti x27 x1 -1862      ====        slti s11, ra, -1862
                                                  30'd    10219    : data = 32'h    016CCB33    ;    //    xor x22 x25 x22      ====        xor s6, s9, s6
                                                  30'd    10220    : data = 32'h    01E020B3    ;    //    slt x1 x0 x30      ====        slt ra, zero, t5
                                                  30'd    10221    : data = 32'h    2F2A7E13    ;    //    andi x28 x20 754      ====        andi t3, s4, 754
                                                  30'd    10222    : data = 32'h    634B2C13    ;    //    slti x24 x22 1588      ====        slti s8, s6, 1588
                                                  30'd    10223    : data = 32'h    0E1A2A37    ;    //    lui x20 57762      ====        lui s4, 57762
                                                  30'd    10224    : data = 32'h    000ED813    ;    //    srli x16 x29 0      ====        srli a6, t4, 0
                                                  30'd    10225    : data = 32'h    C3AEB413    ;    //    sltiu x8 x29 -966      ====        sltiu s0, t4, -966
                                                  30'd    10226    : data = 32'h    0C794893    ;    //    xori x17 x18 199      ====        xori a7, s2, 199
                                                  30'd    10227    : data = 32'h    412857B3    ;    //    sra x15 x16 x18      ====        sra a5, a6, s2
                                                  30'd    10228    : data = 32'h    B6303413    ;    //    sltiu x8 x0 -1181      ====        sltiu s0, zero, -1181
                                                  30'd    10229    : data = 32'h    40D280B3    ;    //    sub x1 x5 x13      ====        sub ra, t0, a3
                                                  30'd    10230    : data = 32'h    00D72CB3    ;    //    slt x25 x14 x13      ====        slt s9, a4, a3
                                                  30'd    10231    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10232    : data = 32'h    B3277E37    ;    //    lui x28 733815      ====        lui t3, 733815
                                                  30'd    10233    : data = 32'h    F3B8E613    ;    //    ori x12 x17 -197      ====        ori a2, a7, -197
                                                  30'd    10234    : data = 32'h    009449B3    ;    //    xor x19 x8 x9      ====        xor s3, s0, s1
                                                  30'd    10235    : data = 32'h    40F0DE93    ;    //    srai x29 x1 15      ====        srai t4, ra, 15
                                                  30'd    10236    : data = 32'h    012AE2B3    ;    //    or x5 x21 x18      ====        or t0, s5, s2
                                                  30'd    10237    : data = 32'h    91D9B813    ;    //    sltiu x16 x19 -1763      ====        sltiu a6, s3, -1763
                                                  30'd    10238    : data = 32'h    E812F613    ;    //    andi x12 x5 -383      ====        andi a2, t0, -383
                                                  30'd    10239    : data = 32'h    00DBFD33    ;    //    and x26 x23 x13      ====        and s10, s7, a3
                                                  30'd    10240    : data = 32'h    00C9DE93    ;    //    srli x29 x19 12      ====        srli t4, s3, 12
                                                  30'd    10241    : data = 32'h    00DD74B3    ;    //    and x9 x26 x13      ====        and s1, s10, a3
                                                  30'd    10242    : data = 32'h    007F5333    ;    //    srl x6 x30 x7      ====        srl t1, t5, t2
                                                  30'd    10243    : data = 32'h    01541A13    ;    //    slli x20 x8 21      ====        slli s4, s0, 21
                                                  30'd    10244    : data = 32'h    00DDD1B3    ;    //    srl x3 x27 x13      ====        srl gp, s11, a3
                                                  30'd    10245    : data = 32'h    41CC5A33    ;    //    sra x20 x24 x28      ====        sra s4, s8, t3
                                                  30'd    10246    : data = 32'h    01EC7833    ;    //    and x16 x24 x30      ====        and a6, s8, t5
                                                  30'd    10247    : data = 32'h    002396B3    ;    //    sll x13 x7 x2      ====        sll a3, t2, sp
                                                  30'd    10248    : data = 32'h    00BB98B3    ;    //    sll x17 x23 x11      ====        sll a7, s7, a1
                                                  30'd    10249    : data = 32'h    8D368713    ;    //    addi x14 x13 -1837      ====        addi a4, a3, -1837
                                                  30'd    10250    : data = 32'h    41125D33    ;    //    sra x26 x4 x17      ====        sra s10, tp, a7
                                                  30'd    10251    : data = 32'h    00B95B93    ;    //    srli x23 x18 11      ====        srli s7, s2, 11
                                                  30'd    10252    : data = 32'h    4A82CF93    ;    //    xori x31 x5 1192      ====        xori t6, t0, 1192
                                                  30'd    10253    : data = 32'h    41065293    ;    //    srai x5 x12 16      ====        srai t0, a2, 16
                                                  30'd    10254    : data = 32'h    00FD8B33    ;    //    add x22 x27 x15      ====        add s6, s11, a5
                                                  30'd    10255    : data = 32'h    00C0B133    ;    //    sltu x2 x1 x12      ====        sltu sp, ra, a2
                                                  30'd    10256    : data = 32'h    04C3C493    ;    //    xori x9 x7 76      ====        xori s1, t2, 76
                                                  30'd    10257    : data = 32'h    47CB5117    ;    //    auipc x2 294069      ====        auipc sp, 294069
                                                  30'd    10258    : data = 32'h    01BF8333    ;    //    add x6 x31 x27      ====        add t1, t6, s11
                                                  30'd    10259    : data = 32'h    C9746B97    ;    //    auipc x23 825158      ====        auipc s7, 825158
                                                  30'd    10260    : data = 32'h    017DE733    ;    //    or x14 x27 x23      ====        or a4, s11, s7
                                                  30'd    10261    : data = 32'h    0160DEB3    ;    //    srl x29 x1 x22      ====        srl t4, ra, s6
                                                  30'd    10262    : data = 32'h    40EF8733    ;    //    sub x14 x31 x14      ====        sub a4, t6, a4
                                                  30'd    10263    : data = 32'h    00EEEA33    ;    //    or x20 x29 x14      ====        or s4, t4, a4
                                                  30'd    10264    : data = 32'h    01000633    ;    //    add x12 x0 x16      ====        add a2, zero, a6
                                                  30'd    10265    : data = 32'h    01DE8FB3    ;    //    add x31 x29 x29      ====        add t6, t4, t4
                                                  30'd    10266    : data = 32'h    0180DCB3    ;    //    srl x25 x1 x24      ====        srl s9, ra, s8
                                                  30'd    10267    : data = 32'h    00C91693    ;    //    slli x13 x18 12      ====        slli a3, s2, 12
                                                  30'd    10268    : data = 32'h    00698EB3    ;    //    add x29 x19 x6      ====        add t4, s3, t1
                                                  30'd    10269    : data = 32'h    015F9DB3    ;    //    sll x27 x31 x21      ====        sll s11, t6, s5
                                                  30'd    10270    : data = 32'h    41310B33    ;    //    sub x22 x2 x19      ====        sub s6, sp, s3
                                                  30'd    10271    : data = 32'h    014A0C33    ;    //    add x24 x20 x20      ====        add s8, s4, s4
                                                  30'd    10272    : data = 32'h    EC89C293    ;    //    xori x5 x19 -312      ====        xori t0, s3, -312
                                                  30'd    10273    : data = 32'h    DD9ACEB7    ;    //    lui x29 907692      ====        lui t4, 907692
                                                  30'd    10274    : data = 32'h    41E3D1B3    ;    //    sra x3 x7 x30      ====        sra gp, t2, t5
                                                  30'd    10275    : data = 32'h    019E7FB3    ;    //    and x31 x28 x25      ====        and t6, t3, s9
                                                  30'd    10276    : data = 32'h    01A07D33    ;    //    and x26 x0 x26      ====        and s10, zero, s10
                                                  30'd    10277    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10278    : data = 32'h    00D488B3    ;    //    add x17 x9 x13      ====        add a7, s1, a3
                                                  30'd    10279    : data = 32'h    40655B13    ;    //    srai x22 x10 6      ====        srai s6, a0, 6
                                                  30'd    10280    : data = 32'h    00BCB133    ;    //    sltu x2 x25 x11      ====        sltu sp, s9, a1
                                                  30'd    10281    : data = 32'h    00DEE7B3    ;    //    or x15 x29 x13      ====        or a5, t4, a3
                                                  30'd    10282    : data = 32'h    48116393    ;    //    ori x7 x2 1153      ====        ori t2, sp, 1153
                                                  30'd    10283    : data = 32'h    00E5E933    ;    //    or x18 x11 x14      ====        or s2, a1, a4
                                                  30'd    10284    : data = 32'h    FF7DE193    ;    //    ori x3 x27 -9      ====        ori gp, s11, -9
                                                  30'd    10285    : data = 32'h    01FD5F93    ;    //    srli x31 x26 31      ====        srli t6, s10, 31
                                                  30'd    10286    : data = 32'h    E7F4A093    ;    //    slti x1 x9 -385      ====        slti ra, s1, -385
                                                  30'd    10287    : data = 32'h    416EDC93    ;    //    srai x25 x29 22      ====        srai s9, t4, 22
                                                  30'd    10288    : data = 32'h    00D580B3    ;    //    add x1 x11 x13      ====        add ra, a1, a3
                                                  30'd    10289    : data = 32'h    01C9AA33    ;    //    slt x20 x19 x28      ====        slt s4, s3, t3
                                                  30'd    10290    : data = 32'h    642C7E37    ;    //    lui x28 410311      ====        lui t3, 410311
                                                  30'd    10291    : data = 32'h    0147AB33    ;    //    slt x22 x15 x20      ====        slt s6, a5, s4
                                                  30'd    10292    : data = 32'h    46D37F93    ;    //    andi x31 x6 1133      ====        andi t6, t1, 1133
                                                  30'd    10293    : data = 32'h    010E2133    ;    //    slt x2 x28 x16      ====        slt sp, t3, a6
                                                  30'd    10294    : data = 32'h    0149D9B3    ;    //    srl x19 x19 x20      ====        srl s3, s3, s4
                                                  30'd    10295    : data = 32'h    90FCC893    ;    //    xori x17 x25 -1777      ====        xori a7, s9, -1777
                                                  30'd    10296    : data = 32'h    22508093    ;    //    addi x1 x1 549      ====        addi ra, ra, 549
                                                  30'd    10297    : data = 32'h    56F06C13    ;    //    ori x24 x0 1391      ====        ori s8, zero, 1391
                                                  30'd    10298    : data = 32'h    59138613    ;    //    addi x12 x7 1425      ====        addi a2, t2, 1425
                                                  30'd    10299    : data = 32'h    00F07EB3    ;    //    and x29 x0 x15      ====        and t4, zero, a5
                                                  30'd    10300    : data = 32'h    40B35113    ;    //    srai x2 x6 11      ====        srai sp, t1, 11
                                                  30'd    10301    : data = 32'h    00F66BB3    ;    //    or x23 x12 x15      ====        or s7, a2, a5
                                                  30'd    10302    : data = 32'h    40C650B3    ;    //    sra x1 x12 x12      ====        sra ra, a2, a2
                                                  30'd    10303    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10304    : data = 32'h    40E35933    ;    //    sra x18 x6 x14      ====        sra s2, t1, a4
                                                  30'd    10305    : data = 32'h    F9322D13    ;    //    slti x26 x4 -109      ====        slti s10, tp, -109
                                                  30'd    10306    : data = 32'h    3CE17013    ;    //    andi x0 x2 974      ====        andi zero, sp, 974
                                                  30'd    10307    : data = 32'h    01EB63B3    ;    //    or x7 x22 x30      ====        or t2, s6, t5
                                                  30'd    10308    : data = 32'h    9AE68E37    ;    //    lui x28 634472      ====        lui t3, 634472
                                                  30'd    10309    : data = 32'h    5A254E13    ;    //    xori x28 x10 1442      ====        xori t3, a0, 1442
                                                  30'd    10310    : data = 32'h    01716FB3    ;    //    or x31 x2 x23      ====        or t6, sp, s7
                                                  30'd    10311    : data = 32'h    41F35D33    ;    //    sra x26 x6 x31      ====        sra s10, t1, t6
                                                  30'd    10312    : data = 32'h    8BEE2597    ;    //    auipc x11 573154      ====        auipc a1, 573154
                                                  30'd    10313    : data = 32'h    411103B3    ;    //    sub x7 x2 x17      ====        sub t2, sp, a7
                                                  30'd    10314    : data = 32'h    89612E13    ;    //    slti x28 x2 -1898      ====        slti t3, sp, -1898
                                                  30'd    10315    : data = 32'h    26E16D13    ;    //    ori x26 x2 622      ====        ori s10, sp, 622
                                                  30'd    10316    : data = 32'h    001707B3    ;    //    add x15 x14 x1      ====        add a5, a4, ra
                                                  30'd    10317    : data = 32'h    000129B3    ;    //    slt x19 x2 x0      ====        slt s3, sp, zero
                                                  30'd    10318    : data = 32'h    41C25133    ;    //    sra x2 x4 x28      ====        sra sp, tp, t3
                                                  30'd    10319    : data = 32'h    01B79933    ;    //    sll x18 x15 x27      ====        sll s2, a5, s11
                                                  30'd    10320    : data = 32'h    8B96CC93    ;    //    xori x25 x13 -1863      ====        xori s9, a3, -1863
                                                  30'd    10321    : data = 32'h    A60B6993    ;    //    ori x19 x22 -1440      ====        ori s3, s6, -1440
                                                  30'd    10322    : data = 32'h    31BC7997    ;    //    auipc x19 203719      ====        auipc s3, 203719
                                                  30'd    10323    : data = 32'h    C378AE93    ;    //    slti x29 x17 -969      ====        slti t4, a7, -969
                                                  30'd    10324    : data = 32'h    0105F0B3    ;    //    and x1 x11 x16      ====        and ra, a1, a6
                                                  30'd    10325    : data = 32'h    858D6493    ;    //    ori x9 x26 -1960      ====        ori s1, s10, -1960
                                                  30'd    10326    : data = 32'h    005BD733    ;    //    srl x14 x23 x5      ====        srl a4, s7, t0
                                                  30'd    10327    : data = 32'h    915B6437    ;    //    lui x8 595382      ====        lui s0, 595382
                                                  30'd    10328    : data = 32'h    01F3DE13    ;    //    srli x28 x7 31      ====        srli t3, t2, 31
                                                  30'd    10329    : data = 32'h    01C0F9B3    ;    //    and x19 x1 x28      ====        and s3, ra, t3
                                                  30'd    10330    : data = 32'h    009B16B3    ;    //    sll x13 x22 x9      ====        sll a3, s6, s1
                                                  30'd    10331    : data = 32'h    00C4A433    ;    //    slt x8 x9 x12      ====        slt s0, s1, a2
                                                  30'd    10332    : data = 32'h    01912E33    ;    //    slt x28 x2 x25      ====        slt t3, sp, s9
                                                  30'd    10333    : data = 32'h    003C7433    ;    //    and x8 x24 x3      ====        and s0, s8, gp
                                                  30'd    10334    : data = 32'h    016B1633    ;    //    sll x12 x22 x22      ====        sll a2, s6, s6
                                                  30'd    10335    : data = 32'h    009EF4B3    ;    //    and x9 x29 x9      ====        and s1, t4, s1
                                                  30'd    10336    : data = 32'h    53023793    ;    //    sltiu x15 x4 1328      ====        sltiu a5, tp, 1328
                                                  30'd    10337    : data = 32'h    00C448B3    ;    //    xor x17 x8 x12      ====        xor a7, s0, a2
                                                  30'd    10338    : data = 32'h    0089A3B3    ;    //    slt x7 x19 x8      ====        slt t2, s3, s0
                                                  30'd    10339    : data = 32'h    01594B33    ;    //    xor x22 x18 x21      ====        xor s6, s2, s5
                                                  30'd    10340    : data = 32'h    00B1BCB3    ;    //    sltu x25 x3 x11      ====        sltu s9, gp, a1
                                                  30'd    10341    : data = 32'h    248EE837    ;    //    lui x16 149742      ====        lui a6, 149742
                                                  30'd    10342    : data = 32'h    41265693    ;    //    srai x13 x12 18      ====        srai a3, a2, 18
                                                  30'd    10343    : data = 32'h    E2F70593    ;    //    addi x11 x14 -465      ====        addi a1, a4, -465
                                                  30'd    10344    : data = 32'h    01871C33    ;    //    sll x24 x14 x24      ====        sll s8, a4, s8
                                                  30'd    10345    : data = 32'h    325F3113    ;    //    sltiu x2 x30 805      ====        sltiu sp, t5, 805
                                                  30'd    10346    : data = 32'h    01D05AB3    ;    //    srl x21 x0 x29      ====        srl s5, zero, t4
                                                  30'd    10347    : data = 32'h    003EDE33    ;    //    srl x28 x29 x3      ====        srl t3, t4, gp
                                                  30'd    10348    : data = 32'h    409300B3    ;    //    sub x1 x6 x9      ====        sub ra, t1, s1
                                                  30'd    10349    : data = 32'h    01502633    ;    //    slt x12 x0 x21      ====        slt a2, zero, s5
                                                  30'd    10350    : data = 32'h    16FF23B7    ;    //    lui x7 94194      ====        lui t2, 94194
                                                  30'd    10351    : data = 32'h    0189ED33    ;    //    or x26 x19 x24      ====        or s10, s3, s8
                                                  30'd    10352    : data = 32'h    01435433    ;    //    srl x8 x6 x20      ====        srl s0, t1, s4
                                                  30'd    10353    : data = 32'h    00D380B3    ;    //    add x1 x7 x13      ====        add ra, t2, a3
                                                  30'd    10354    : data = 32'h    F2C6A913    ;    //    slti x18 x13 -212      ====        slti s2, a3, -212
                                                  30'd    10355    : data = 32'h    017511B3    ;    //    sll x3 x10 x23      ====        sll gp, a0, s7
                                                  30'd    10356    : data = 32'h    01BDBBB3    ;    //    sltu x23 x27 x27      ====        sltu s7, s11, s11
                                                  30'd    10357    : data = 32'h    0B0D6593    ;    //    ori x11 x26 176      ====        ori a1, s10, 176
                                                  30'd    10358    : data = 32'h    C0AEE593    ;    //    ori x11 x29 -1014      ====        ori a1, t4, -1014
                                                  30'd    10359    : data = 32'h    A672AB93    ;    //    slti x23 x5 -1433      ====        slti s7, t0, -1433
                                                  30'd    10360    : data = 32'h    0079B033    ;    //    sltu x0 x19 x7      ====        sltu zero, s3, t2
                                                  30'd    10361    : data = 32'h    0BB76C93    ;    //    ori x25 x14 187      ====        ori s9, a4, 187
                                                  30'd    10362    : data = 32'h    0017E5B3    ;    //    or x11 x15 x1      ====        or a1, a5, ra
                                                  30'd    10363    : data = 32'h    015C6B33    ;    //    or x22 x24 x21      ====        or s6, s8, s5
                                                  30'd    10364    : data = 32'h    0029D993    ;    //    srli x19 x19 2      ====        srli s3, s3, 2
                                                  30'd    10365    : data = 32'h    41A753B3    ;    //    sra x7 x14 x26      ====        sra t2, a4, s10
                                                  30'd    10366    : data = 32'h    00012FB3    ;    //    slt x31 x2 x0      ====        slt t6, sp, zero
                                                  30'd    10367    : data = 32'h    01F895B3    ;    //    sll x11 x17 x31      ====        sll a1, a7, t6
                                                  30'd    10368    : data = 32'h    FB55E893    ;    //    ori x17 x11 -75      ====        ori a7, a1, -75
                                                  30'd    10369    : data = 32'h    012A0333    ;    //    add x6 x20 x18      ====        add t1, s4, s2
                                                  30'd    10370    : data = 32'h    40FF01B3    ;    //    sub x3 x30 x15      ====        sub gp, t5, a5
                                                  30'd    10371    : data = 32'h    E397FA13    ;    //    andi x20 x15 -455      ====        andi s4, a5, -455
                                                  30'd    10372    : data = 32'h    76767093    ;    //    andi x1 x12 1895      ====        andi ra, a2, 1895
                                                  30'd    10373    : data = 32'h    40A0D893    ;    //    srai x17 x1 10      ====        srai a7, ra, 10
                                                  30'd    10374    : data = 32'h    00DA9D33    ;    //    sll x26 x21 x13      ====        sll s10, s5, a3
                                                  30'd    10375    : data = 32'h    00889293    ;    //    slli x5 x17 8      ====        slli t0, a7, 8
                                                  30'd    10376    : data = 32'h    01B25EB3    ;    //    srl x29 x4 x27      ====        srl t4, tp, s11
                                                  30'd    10377    : data = 32'h    011AD4B3    ;    //    srl x9 x21 x17      ====        srl s1, s5, a7
                                                  30'd    10378    : data = 32'h    00A487B3    ;    //    add x15 x9 x10      ====        add a5, s1, a0
                                                  30'd    10379    : data = 32'h    4035D193    ;    //    srai x3 x11 3      ====        srai gp, a1, 3
                                                  30'd    10380    : data = 32'h    41685833    ;    //    sra x16 x16 x22      ====        sra a6, a6, s6
                                                  30'd    10381    : data = 32'h    01DF8E33    ;    //    add x28 x31 x29      ====        add t3, t6, t4
                                                  30'd    10382    : data = 32'h    01008833    ;    //    add x16 x1 x16      ====        add a6, ra, a6
                                                  30'd    10383    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10384    : data = 32'h    0038F833    ;    //    and x16 x17 x3      ====        and a6, a7, gp
                                                  30'd    10385    : data = 32'h    00D97FB3    ;    //    and x31 x18 x13      ====        and t6, s2, a3
                                                  30'd    10386    : data = 32'h    009AB033    ;    //    sltu x0 x21 x9      ====        sltu zero, s5, s1
                                                  30'd    10387    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10388    : data = 32'h    00B88B33    ;    //    add x22 x17 x11      ====        add s6, a7, a1
                                                  30'd    10389    : data = 32'h    005AE933    ;    //    or x18 x21 x5      ====        or s2, s5, t0
                                                  30'd    10390    : data = 32'h    373DB613    ;    //    sltiu x12 x27 883      ====        sltiu a2, s11, 883
                                                  30'd    10391    : data = 32'h    0195C433    ;    //    xor x8 x11 x25      ====        xor s0, a1, s9
                                                  30'd    10392    : data = 32'h    410D0833    ;    //    sub x16 x26 x16      ====        sub a6, s10, a6
                                                  30'd    10393    : data = 32'h    019258B3    ;    //    srl x17 x4 x25      ====        srl a7, tp, s9
                                                  30'd    10394    : data = 32'h    0FFA2293    ;    //    slti x5 x20 255      ====        slti t0, s4, 255
                                                  30'd    10395    : data = 32'h    009D8B33    ;    //    add x22 x27 x9      ====        add s6, s11, s1
                                                  30'd    10396    : data = 32'h    01357D33    ;    //    and x26 x10 x19      ====        and s10, a0, s3
                                                  30'd    10397    : data = 32'h    01725CB3    ;    //    srl x25 x4 x23      ====        srl s9, tp, s7
                                                  30'd    10398    : data = 32'h    01AD9133    ;    //    sll x2 x27 x26      ====        sll sp, s11, s10
                                                  30'd    10399    : data = 32'h    16ABF593    ;    //    andi x11 x23 362      ====        andi a1, s7, 362
                                                  30'd    10400    : data = 32'h    01D2EBB3    ;    //    or x23 x5 x29      ====        or s7, t0, t4
                                                  30'd    10401    : data = 32'h    017345B3    ;    //    xor x11 x6 x23      ====        xor a1, t1, s7
                                                  30'd    10402    : data = 32'h    FFF00D93    ;    //    addi x27 x0 -1      ====        li s11, 0xffffffff #start riscv_int_numeric_corner_stream_30
                                                  30'd    10403    : data = 32'h    B8631C37    ;    //    lui x24 755249      ====        li s8, 0xb8630f0a
                                                  30'd    10404    : data = 32'h    F0AC0C13    ;    //    addi x24 x24 -246      ====        li s8, 0xb8630f0a
                                                  30'd    10405    : data = 32'h    83D24BB7    ;    //    lui x23 539940      ====        li s7, 0x83d23a08
                                                  30'd    10406    : data = 32'h    A08B8B93    ;    //    addi x23 x23 -1528      ====        li s7, 0x83d23a08
                                                  30'd    10407    : data = 32'h    00000693    ;    //    addi x13 x0 0      ====        li a3, 0x0
                                                  30'd    10408    : data = 32'h    80000FB7    ;    //    lui x31 524288      ====        li t6, 0x80000000
                                                  30'd    10409    : data = 32'h    000F8F93    ;    //    addi x31 x31 0      ====        li t6, 0x80000000
                                                  30'd    10410    : data = 32'h    800002B7    ;    //    lui x5 524288      ====        li t0, 0x80000000
                                                  30'd    10411    : data = 32'h    00028293    ;    //    addi x5 x5 0      ====        li t0, 0x80000000
                                                  30'd    10412    : data = 32'h    00000493    ;    //    addi x9 x0 0      ====        li s1, 0x0
                                                  30'd    10413    : data = 32'h    E1781E37    ;    //    lui x28 923521      ====        li t3, 0xe17814c6
                                                  30'd    10414    : data = 32'h    4C6E0E13    ;    //    addi x28 x28 1222      ====        li t3, 0xe17814c6
                                                  30'd    10415    : data = 32'h    00000813    ;    //    addi x16 x0 0      ====        li a6, 0x0
                                                  30'd    10416    : data = 32'h    00000593    ;    //    addi x11 x0 0      ====        li a1, 0x0
                                                  30'd    10417    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10418    : data = 32'h    D26B7817    ;    //    auipc x16 861879      ====        auipc a6, 861879
                                                  30'd    10419    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10420    : data = 32'h    00BC04B3    ;    //    add x9 x24 x11      ====        add s1, s8, a1
                                                  30'd    10421    : data = 32'h    B5D75D97    ;    //    auipc x27 744821      ====        auipc s11, 744821
                                                  30'd    10422    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10423    : data = 32'h    40DC06B3    ;    //    sub x13 x24 x13      ====        sub a3, s8, a3
                                                  30'd    10424    : data = 32'h    787C1817    ;    //    auipc x16 493505      ====        auipc a6, 493505
                                                  30'd    10425    : data = 32'h    7892F497    ;    //    auipc x9 493871      ====        auipc s1, 493871
                                                  30'd    10426    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10427    : data = 32'h    41CD85B3    ;    //    sub x11 x27 x28      ====        sub a1, s11, t3
                                                  30'd    10428    : data = 32'h    90FDC817    ;    //    auipc x16 593884      ====        auipc a6, 593884
                                                  30'd    10429    : data = 32'h    814AF5B7    ;    //    lui x11 529583      ====        lui a1, 529583
                                                  30'd    10430    : data = 32'h    01F482B3    ;    //    add x5 x9 x31      ====        add t0, s1, t6
                                                  30'd    10431    : data = 32'h    8032F6B7    ;    //    lui x13 525103      ====        lui a3, 525103
                                                  30'd    10432    : data = 32'h    00BD8FB3    ;    //    add x31 x27 x11      ====        add t6, s11, a1
                                                  30'd    10433    : data = 32'h    410D8E33    ;    //    sub x28 x27 x16      ====        sub t3, s11, a6
                                                  30'd    10434    : data = 32'h    00DC05B3    ;    //    add x11 x24 x13      ====        add a1, s8, a3
                                                  30'd    10435    : data = 32'h    138C0813    ;    //    addi x16 x24 312      ====        addi a6, s8, 312
                                                  30'd    10436    : data = 32'h    BEE28493    ;    //    addi x9 x5 -1042      ====        addi s1, t0, -1042
                                                  30'd    10437    : data = 32'h    017D86B3    ;    //    add x13 x27 x23      ====        add a3, s11, s7
                                                  30'd    10438    : data = 32'h    41880C33    ;    //    sub x24 x16 x24      ====        sub s8, a6, s8
                                                  30'd    10439    : data = 32'h    009B8FB3    ;    //    add x31 x23 x9      ====        add t6, s7, s1
                                                  30'd    10440    : data = 32'h    DFCB74B7    ;    //    lui x9 916663      ====        lui s1, 916663
                                                  30'd    10441    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10442    : data = 32'h    21A1C4B7    ;    //    lui x9 137756      ====        lui s1, 137756
                                                  30'd    10443    : data = 32'h    410CEC37    ;    //    lui x24 266446      ====        lui s8, 266446
                                                  30'd    10444    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10445    : data = 32'h    3B4010EF    ;    //    jal x1 5044      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_30
                                                  30'd    10446    : data = 32'h    DC42FD93    ;    //    andi x27 x5 -572      ====        andi s11, t0, -572
                                                  30'd    10447    : data = 32'h    00ABD7B3    ;    //    srl x15 x23 x10      ====        srl a5, s7, a0
                                                  30'd    10448    : data = 32'h    C08B6313    ;    //    ori x6 x22 -1016      ====        ori t1, s6, -1016
                                                  30'd    10449    : data = 32'h    0173F433    ;    //    and x8 x7 x23      ====        and s0, t2, s7
                                                  30'd    10450    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10451    : data = 32'h    4157D4B3    ;    //    sra x9 x15 x21      ====        sra s1, a5, s5
                                                  30'd    10452    : data = 32'h    00DC34B3    ;    //    sltu x9 x24 x13      ====        sltu s1, s8, a3
                                                  30'd    10453    : data = 32'h    0147DEB3    ;    //    srl x29 x15 x20      ====        srl t4, a5, s4
                                                  30'd    10454    : data = 32'h    CD3F7613    ;    //    andi x12 x30 -813      ====        andi a2, t5, -813
                                                  30'd    10455    : data = 32'h    AD007813    ;    //    andi x16 x0 -1328      ====        andi a6, zero, -1328
                                                  30'd    10456    : data = 32'h    0161D2B3    ;    //    srl x5 x3 x22      ====        srl t0, gp, s6
                                                  30'd    10457    : data = 32'h    00154733    ;    //    xor x14 x10 x1      ====        xor a4, a0, ra
                                                  30'd    10458    : data = 32'h    00F26B33    ;    //    or x22 x4 x15      ====        or s6, tp, a5
                                                  30'd    10459    : data = 32'h    7ED9FCB7    ;    //    lui x25 519583      ====        lui s9, 519583
                                                  30'd    10460    : data = 32'h    019A1133    ;    //    sll x2 x20 x25      ====        sll sp, s4, s9
                                                  30'd    10461    : data = 32'h    4C163EB7    ;    //    lui x29 311651      ====        lui t4, 311651
                                                  30'd    10462    : data = 32'h    00D0E7B3    ;    //    or x15 x1 x13      ====        or a5, ra, a3
                                                  30'd    10463    : data = 32'h    000A6AB3    ;    //    or x21 x20 x0      ====        or s5, s4, zero
                                                  30'd    10464    : data = 32'h    01FB9313    ;    //    slli x6 x23 31      ====        slli t1, s7, 31
                                                  30'd    10465    : data = 32'h    FE770893    ;    //    addi x17 x14 -25      ====        addi a7, a4, -25
                                                  30'd    10466    : data = 32'h    DDB8C713    ;    //    xori x14 x17 -549      ====        xori a4, a7, -549
                                                  30'd    10467    : data = 32'h    00935193    ;    //    srli x3 x6 9      ====        srli gp, t1, 9
                                                  30'd    10468    : data = 32'h    ABB42713    ;    //    slti x14 x8 -1349      ====        slti a4, s0, -1349
                                                  30'd    10469    : data = 32'h    CE21EC13    ;    //    ori x24 x3 -798      ====        ori s8, gp, -798
                                                  30'd    10470    : data = 32'h    243AC613    ;    //    xori x12 x21 579      ====        xori a2, s5, 579
                                                  30'd    10471    : data = 32'h    01EBBAB3    ;    //    sltu x21 x23 x30      ====        sltu s5, s7, t5
                                                  30'd    10472    : data = 32'h    C7F82997    ;    //    auipc x19 819074      ====        auipc s3, 819074
                                                  30'd    10473    : data = 32'h    EB437D93    ;    //    andi x27 x6 -332      ====        andi s11, t1, -332
                                                  30'd    10474    : data = 32'h    001E1893    ;    //    slli x17 x28 1      ====        slli a7, t3, 1
                                                  30'd    10475    : data = 32'h    2BBA4937    ;    //    lui x18 179108      ====        lui s2, 179108
                                                  30'd    10476    : data = 32'h    004DD013    ;    //    srli x0 x27 4      ====        srli zero, s11, 4
                                                  30'd    10477    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10478    : data = 32'h    01B4ED33    ;    //    or x26 x9 x27      ====        or s10, s1, s11
                                                  30'd    10479    : data = 32'h    01BC1B13    ;    //    slli x22 x24 27      ====        slli s6, s8, 27
                                                  30'd    10480    : data = 32'h    00314433    ;    //    xor x8 x2 x3      ====        xor s0, sp, gp
                                                  30'd    10481    : data = 32'h    8142F713    ;    //    andi x14 x5 -2028      ====        andi a4, t0, -2028
                                                  30'd    10482    : data = 32'h    004E5733    ;    //    srl x14 x28 x4      ====        srl a4, t3, tp
                                                  30'd    10483    : data = 32'h    01C26733    ;    //    or x14 x4 x28      ====        or a4, tp, t3
                                                  30'd    10484    : data = 32'h    00E878B3    ;    //    and x17 x16 x14      ====        and a7, a6, a4
                                                  30'd    10485    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10486    : data = 32'h    40FC0DB3    ;    //    sub x27 x24 x15      ====        sub s11, s8, a5
                                                  30'd    10487    : data = 32'h    01D2D393    ;    //    srli x7 x5 29      ====        srli t2, t0, 29
                                                  30'd    10488    : data = 32'h    01A72DB3    ;    //    slt x27 x14 x26      ====        slt s11, a4, s10
                                                  30'd    10489    : data = 32'h    00F29D13    ;    //    slli x26 x5 15      ====        slli s10, t0, 15
                                                  30'd    10490    : data = 32'h    00BE5413    ;    //    srli x8 x28 11      ====        srli s0, t3, 11
                                                  30'd    10491    : data = 32'h    01A4BB33    ;    //    sltu x22 x9 x26      ====        sltu s6, s1, s10
                                                  30'd    10492    : data = 32'h    ACEF0D13    ;    //    addi x26 x30 -1330      ====        addi s10, t5, -1330
                                                  30'd    10493    : data = 32'h    C33BA813    ;    //    slti x16 x23 -973      ====        slti a6, s7, -973
                                                  30'd    10494    : data = 32'h    005B51B3    ;    //    srl x3 x22 x5      ====        srl gp, s6, t0
                                                  30'd    10495    : data = 32'h    41915693    ;    //    srai x13 x2 25      ====        srai a3, sp, 25
                                                  30'd    10496    : data = 32'h    01B792B3    ;    //    sll x5 x15 x27      ====        sll t0, a5, s11
                                                  30'd    10497    : data = 32'h    52563017    ;    //    auipc x0 337251      ====        auipc zero, 337251
                                                  30'd    10498    : data = 32'h    01D90733    ;    //    add x14 x18 x29      ====        add a4, s2, t4
                                                  30'd    10499    : data = 32'h    907FF093    ;    //    andi x1 x31 -1785      ====        andi ra, t6, -1785
                                                  30'd    10500    : data = 32'h    003AA933    ;    //    slt x18 x21 x3      ====        slt s2, s5, gp
                                                  30'd    10501    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10502    : data = 32'h    40370DB3    ;    //    sub x27 x14 x3      ====        sub s11, a4, gp
                                                  30'd    10503    : data = 32'h    6F155F97    ;    //    auipc x31 454997      ====        auipc t6, 454997
                                                  30'd    10504    : data = 32'h    41A5D413    ;    //    srai x8 x11 26      ====        srai s0, a1, 26
                                                  30'd    10505    : data = 32'h    D893FB93    ;    //    andi x23 x7 -631      ====        andi s7, t2, -631
                                                  30'd    10506    : data = 32'h    838798B7    ;    //    lui x17 538745      ====        lui a7, 538745
                                                  30'd    10507    : data = 32'h    99BC3B97    ;    //    auipc x23 629699      ====        auipc s7, 629699
                                                  30'd    10508    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10509    : data = 32'h    41ADD913    ;    //    srai x18 x27 26      ====        srai s2, s11, 26
                                                  30'd    10510    : data = 32'h    00E5B1B3    ;    //    sltu x3 x11 x14      ====        sltu gp, a1, a4
                                                  30'd    10511    : data = 32'h    00DF0BB3    ;    //    add x23 x30 x13      ====        add s7, t5, a3
                                                  30'd    10512    : data = 32'h    1A3B4D97    ;    //    auipc x27 107444      ====        auipc s11, 107444
                                                  30'd    10513    : data = 32'h    05D76A13    ;    //    ori x20 x14 93      ====        ori s4, a4, 93
                                                  30'd    10514    : data = 32'h    001B5833    ;    //    srl x16 x22 x1      ====        srl a6, s6, ra
                                                  30'd    10515    : data = 32'h    D0DCAA93    ;    //    slti x21 x25 -755      ====        slti s5, s9, -755
                                                  30'd    10516    : data = 32'h    B126A493    ;    //    slti x9 x13 -1262      ====        slti s1, a3, -1262
                                                  30'd    10517    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10518    : data = 32'h    C895BE13    ;    //    sltiu x28 x11 -887      ====        sltiu t3, a1, -887
                                                  30'd    10519    : data = 32'h    00768933    ;    //    add x18 x13 x7      ====        add s2, a3, t2
                                                  30'd    10520    : data = 32'h    00E25F93    ;    //    srli x31 x4 14      ====        srli t6, tp, 14
                                                  30'd    10521    : data = 32'h    424CC913    ;    //    xori x18 x25 1060      ====        xori s2, s9, 1060
                                                  30'd    10522    : data = 32'h    01B749B3    ;    //    xor x19 x14 x27      ====        xor s3, a4, s11
                                                  30'd    10523    : data = 32'h    FDD1C893    ;    //    xori x17 x3 -35      ====        xori a7, gp, -35
                                                  30'd    10524    : data = 32'h    E0E82113    ;    //    slti x2 x16 -498      ====        slti sp, a6, -498
                                                  30'd    10525    : data = 32'h    01FB8033    ;    //    add x0 x23 x31      ====        add zero, s7, t6
                                                  30'd    10526    : data = 32'h    C3B91E37    ;    //    lui x28 801681      ====        li t3, 0xc3b90df8 #start riscv_int_numeric_corner_stream_28
                                                  30'd    10527    : data = 32'h    DF8E0E13    ;    //    addi x28 x28 -520      ====        li t3, 0xc3b90df8 #start riscv_int_numeric_corner_stream_28
                                                  30'd    10528    : data = 32'h    6FD838B7    ;    //    lui x17 458115      ====        li a7, 0x6fd82f9b
                                                  30'd    10529    : data = 32'h    F9B88893    ;    //    addi x17 x17 -101      ====        li a7, 0x6fd82f9b
                                                  30'd    10530    : data = 32'h    00000193    ;    //    addi x3 x0 0      ====        li gp, 0x0
                                                  30'd    10531    : data = 32'h    00000093    ;    //    addi x1 x0 0      ====        li ra, 0x0
                                                  30'd    10532    : data = 32'h    C0E697B7    ;    //    lui x15 790121      ====        li a5, 0xc0e697f6
                                                  30'd    10533    : data = 32'h    7F678793    ;    //    addi x15 x15 2038      ====        li a5, 0xc0e697f6
                                                  30'd    10534    : data = 32'h    00000713    ;    //    addi x14 x0 0      ====        li a4, 0x0
                                                  30'd    10535    : data = 32'h    00000D93    ;    //    addi x27 x0 0      ====        li s11, 0x0
                                                  30'd    10536    : data = 32'h    BC273C37    ;    //    lui x24 770675      ====        li s8, 0xbc2730f7
                                                  30'd    10537    : data = 32'h    0F7C0C13    ;    //    addi x24 x24 247      ====        li s8, 0xbc2730f7
                                                  30'd    10538    : data = 32'h    865C06B7    ;    //    lui x13 550336      ====        li a3, 0x865bfe0d
                                                  30'd    10539    : data = 32'h    E0D68693    ;    //    addi x13 x13 -499      ====        li a3, 0x865bfe0d
                                                  30'd    10540    : data = 32'h    DB627D37    ;    //    lui x26 898599      ====        li s10, 0xdb626fd2
                                                  30'd    10541    : data = 32'h    FD2D0D13    ;    //    addi x26 x26 -46      ====        li s10, 0xdb626fd2
                                                  30'd    10542    : data = 32'h    E6E32C37    ;    //    lui x24 945714      ====        lui s8, 945714
                                                  30'd    10543    : data = 32'h    24D88D13    ;    //    addi x26 x17 589      ====        addi s10, a7, 589
                                                  30'd    10544    : data = 32'h    E0BD5897    ;    //    auipc x17 920533      ====        auipc a7, 920533
                                                  30'd    10545    : data = 32'h    43268D93    ;    //    addi x27 x13 1074      ====        addi s11, a3, 1074
                                                  30'd    10546    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10547    : data = 32'h    41A881B3    ;    //    sub x3 x17 x26      ====        sub gp, a7, s10
                                                  30'd    10548    : data = 32'h    95BCA6B7    ;    //    lui x13 613322      ====        lui a3, 613322
                                                  30'd    10549    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10550    : data = 32'h    00DD87B3    ;    //    add x15 x27 x13      ====        add a5, s11, a3
                                                  30'd    10551    : data = 32'h    BF580D37    ;    //    lui x26 783744      ====        lui s10, 783744
                                                  30'd    10552    : data = 32'h    4B252097    ;    //    auipc x1 307794      ====        auipc ra, 307794
                                                  30'd    10553    : data = 32'h    00F70E33    ;    //    add x28 x14 x15      ====        add t3, a4, a5
                                                  30'd    10554    : data = 32'h    6B325D37    ;    //    lui x26 439077      ====        lui s10, 439077
                                                  30'd    10555    : data = 32'h    BC8D0093    ;    //    addi x1 x26 -1080      ====        addi ra, s10, -1080
                                                  30'd    10556    : data = 32'h    401E00B3    ;    //    sub x1 x28 x1      ====        sub ra, t3, ra
                                                  30'd    10557    : data = 32'h    E55A6097    ;    //    auipc x1 939430      ====        auipc ra, 939430
                                                  30'd    10558    : data = 32'h    81A80697    ;    //    auipc x13 531072      ====        auipc a3, 531072
                                                  30'd    10559    : data = 32'h    AE7858B7    ;    //    lui x17 714629      ====        lui a7, 714629
                                                  30'd    10560    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10561    : data = 32'h    98B18193    ;    //    addi x3 x3 -1653      ====        addi gp, gp, -1653
                                                  30'd    10562    : data = 32'h    B82240B7    ;    //    lui x1 754212      ====        lui ra, 754212
                                                  30'd    10563    : data = 32'h    E53A66B7    ;    //    lui x13 938918      ====        lui a3, 938918
                                                  30'd    10564    : data = 32'h    E84B78B7    ;    //    lui x17 951479      ====        lui a7, 951479
                                                  30'd    10565    : data = 32'h    40F788B3    ;    //    sub x17 x15 x15      ====        sub a7, a5, a5
                                                  30'd    10566    : data = 32'h    1D0010EF    ;    //    jal x1 4560      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_28
                                                  30'd    10567    : data = 32'h    00315C33    ;    //    srl x24 x2 x3      ====        srl s8, sp, gp
                                                  30'd    10568    : data = 32'h    01FE5D33    ;    //    srl x26 x28 x31      ====        srl s10, t3, t6
                                                  30'd    10569    : data = 32'h    0100FEB3    ;    //    and x29 x1 x16      ====        and t4, ra, a6
                                                  30'd    10570    : data = 32'h    007D2DB3    ;    //    slt x27 x26 x7      ====        slt s11, s10, t2
                                                  30'd    10571    : data = 32'h    3DF88393    ;    //    addi x7 x17 991      ====        addi t2, a7, 991
                                                  30'd    10572    : data = 32'h    0181F6B3    ;    //    and x13 x3 x24      ====        and a3, gp, s8
                                                  30'd    10573    : data = 32'h    5A2E4113    ;    //    xori x2 x28 1442      ====        xori sp, t3, 1442
                                                  30'd    10574    : data = 32'h    01A18B33    ;    //    add x22 x3 x26      ====        add s6, gp, s10
                                                  30'd    10575    : data = 32'h    00DE8133    ;    //    add x2 x29 x13      ====        add sp, t4, a3
                                                  30'd    10576    : data = 32'h    2D040437    ;    //    lui x8 184384      ====        lui s0, 184384
                                                  30'd    10577    : data = 32'h    411304B3    ;    //    sub x9 x6 x17      ====        sub s1, t1, a7
                                                  30'd    10578    : data = 32'h    0072D8B3    ;    //    srl x17 x5 x7      ====        srl a7, t0, t2
                                                  30'd    10579    : data = 32'h    2E684993    ;    //    xori x19 x16 742      ====        xori s3, a6, 742
                                                  30'd    10580    : data = 32'h    402CD993    ;    //    srai x19 x25 2      ====        srai s3, s9, 2
                                                  30'd    10581    : data = 32'h    96465617    ;    //    auipc x12 615525      ====        auipc a2, 615525
                                                  30'd    10582    : data = 32'h    15A43393    ;    //    sltiu x7 x8 346      ====        sltiu t2, s0, 346
                                                  30'd    10583    : data = 32'h    004100B3    ;    //    add x1 x2 x4      ====        add ra, sp, tp
                                                  30'd    10584    : data = 32'h    932E2E93    ;    //    slti x29 x28 -1742      ====        slti t4, t3, -1742
                                                  30'd    10585    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10586    : data = 32'h    20A6BC13    ;    //    sltiu x24 x13 522      ====        sltiu s8, a3, 522
                                                  30'd    10587    : data = 32'h    00187E33    ;    //    and x28 x16 x1      ====        and t3, a6, ra
                                                  30'd    10588    : data = 32'h    009D0133    ;    //    add x2 x26 x9      ====        add sp, s10, s1
                                                  30'd    10589    : data = 32'h    01533E33    ;    //    sltu x28 x6 x21      ====        sltu t3, t1, s5
                                                  30'd    10590    : data = 32'h    00A117B3    ;    //    sll x15 x2 x10      ====        sll a5, sp, a0
                                                  30'd    10591    : data = 32'h    4026D6B3    ;    //    sra x13 x13 x2      ====        sra a3, a3, sp
                                                  30'd    10592    : data = 32'h    DAD3F793    ;    //    andi x15 x7 -595      ====        andi a5, t2, -595
                                                  30'd    10593    : data = 32'h    4003D0B3    ;    //    sra x1 x7 x0      ====        sra ra, t2, zero
                                                  30'd    10594    : data = 32'h    58B56A13    ;    //    ori x20 x10 1419      ====        ori s4, a0, 1419
                                                  30'd    10595    : data = 32'h    D724AA93    ;    //    slti x21 x9 -654      ====        slti s5, s1, -654
                                                  30'd    10596    : data = 32'h    0022D0B3    ;    //    srl x1 x5 x2      ====        srl ra, t0, sp
                                                  30'd    10597    : data = 32'h    012C5FB3    ;    //    srl x31 x24 x18      ====        srl t6, s8, s2
                                                  30'd    10598    : data = 32'h    01F80C33    ;    //    add x24 x16 x31      ====        add s8, a6, t6
                                                  30'd    10599    : data = 32'h    A1384A13    ;    //    xori x20 x16 -1517      ====        xori s4, a6, -1517
                                                  30'd    10600    : data = 32'h    00C19B93    ;    //    slli x23 x3 12      ====        slli s7, gp, 12
                                                  30'd    10601    : data = 32'h    6AA58993    ;    //    addi x19 x11 1706      ====        addi s3, a1, 1706
                                                  30'd    10602    : data = 32'h    00F5AA33    ;    //    slt x20 x11 x15      ====        slt s4, a1, a5
                                                  30'd    10603    : data = 32'h    41C90A33    ;    //    sub x20 x18 x28      ====        sub s4, s2, t3
                                                  30'd    10604    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10605    : data = 32'h    58868193    ;    //    addi x3 x13 1416      ====        addi gp, a3, 1416
                                                  30'd    10606    : data = 32'h    01D90DB3    ;    //    add x27 x18 x29      ====        add s11, s2, t4
                                                  30'd    10607    : data = 32'h    BAB2BD93    ;    //    sltiu x27 x5 -1109      ====        sltiu s11, t0, -1109
                                                  30'd    10608    : data = 32'h    8CF90C93    ;    //    addi x25 x18 -1841      ====        addi s9, s2, -1841
                                                  30'd    10609    : data = 32'h    A5E23693    ;    //    sltiu x13 x4 -1442      ====        sltiu a3, tp, -1442
                                                  30'd    10610    : data = 32'h    01EAD333    ;    //    srl x6 x21 x30      ====        srl t1, s5, t5
                                                  30'd    10611    : data = 32'h    00889693    ;    //    slli x13 x17 8      ====        slli a3, a7, 8
                                                  30'd    10612    : data = 32'h    00A25093    ;    //    srli x1 x4 10      ====        srli ra, tp, 10
                                                  30'd    10613    : data = 32'h    00105433    ;    //    srl x8 x0 x1      ====        srl s0, zero, ra
                                                  30'd    10614    : data = 32'h    07FA4413    ;    //    xori x8 x20 127      ====        xori s0, s4, 127
                                                  30'd    10615    : data = 32'h    41F2D793    ;    //    srai x15 x5 31      ====        srai a5, t0, 31
                                                  30'd    10616    : data = 32'h    016554B3    ;    //    srl x9 x10 x22      ====        srl s1, a0, s6
                                                  30'd    10617    : data = 32'h    00514FB3    ;    //    xor x31 x2 x5      ====        xor t6, sp, t0
                                                  30'd    10618    : data = 32'h    06258A37    ;    //    lui x20 25176      ====        lui s4, 25176
                                                  30'd    10619    : data = 32'h    00870833    ;    //    add x16 x14 x8      ====        add a6, a4, s0
                                                  30'd    10620    : data = 32'h    01E09593    ;    //    slli x11 x1 30      ====        slli a1, ra, 30
                                                  30'd    10621    : data = 32'h    00DB37B3    ;    //    sltu x15 x22 x13      ====        sltu a5, s6, a3
                                                  30'd    10622    : data = 32'h    47A7FF97    ;    //    auipc x31 293503      ====        auipc t6, 293503
                                                  30'd    10623    : data = 32'h    01A48AB3    ;    //    add x21 x9 x26      ====        add s5, s1, s10
                                                  30'd    10624    : data = 32'h    36DFE893    ;    //    ori x17 x31 877      ====        ori a7, t6, 877
                                                  30'd    10625    : data = 32'h    0035D2B3    ;    //    srl x5 x11 x3      ====        srl t0, a1, gp
                                                  30'd    10626    : data = 32'h    14850A13    ;    //    addi x20 x10 328      ====        addi s4, a0, 328
                                                  30'd    10627    : data = 32'h    4190D1B3    ;    //    sra x3 x1 x25      ====        sra gp, ra, s9
                                                  30'd    10628    : data = 32'h    016E9B33    ;    //    sll x22 x29 x22      ====        sll s6, t4, s6
                                                  30'd    10629    : data = 32'h    41870733    ;    //    sub x14 x14 x24      ====        sub a4, a4, s8
                                                  30'd    10630    : data = 32'h    14013D17    ;    //    auipc x26 81939      ====        auipc s10, 81939
                                                  30'd    10631    : data = 32'h    00EDD713    ;    //    srli x14 x27 14      ====        srli a4, s11, 14
                                                  30'd    10632    : data = 32'h    A111BB13    ;    //    sltiu x22 x3 -1519      ====        sltiu s6, gp, -1519
                                                  30'd    10633    : data = 32'h    004E2D33    ;    //    slt x26 x28 x4      ====        slt s10, t3, tp
                                                  30'd    10634    : data = 32'h    B5657493    ;    //    andi x9 x10 -1194      ====        andi s1, a0, -1194
                                                  30'd    10635    : data = 32'h    018C33B3    ;    //    sltu x7 x24 x24      ====        sltu t2, s8, s8
                                                  30'd    10636    : data = 32'h    165B0913    ;    //    addi x18 x22 357      ====        addi s2, s6, 357
                                                  30'd    10637    : data = 32'h    4E74E493    ;    //    ori x9 x9 1255      ====        ori s1, s1, 1255
                                                  30'd    10638    : data = 32'h    406F0133    ;    //    sub x2 x30 x6      ====        sub sp, t5, t1
                                                  30'd    10639    : data = 32'h    98A3EB13    ;    //    ori x22 x7 -1654      ====        ori s6, t2, -1654
                                                  30'd    10640    : data = 32'h    008D1E33    ;    //    sll x28 x26 x8      ====        sll t3, s10, s0
                                                  30'd    10641    : data = 32'h    000F7133    ;    //    and x2 x30 x0      ====        and sp, t5, zero
                                                  30'd    10642    : data = 32'h    29E67013    ;    //    andi x0 x12 670      ====        andi zero, a2, 670
                                                  30'd    10643    : data = 32'h    409A83B3    ;    //    sub x7 x21 x9      ====        sub t2, s5, s1
                                                  30'd    10644    : data = 32'h    00C2C433    ;    //    xor x8 x5 x12      ====        xor s0, t0, a2
                                                  30'd    10645    : data = 32'h    007721B3    ;    //    slt x3 x14 x7      ====        slt gp, a4, t2
                                                  30'd    10646    : data = 32'h    0048B033    ;    //    sltu x0 x17 x4      ====        sltu zero, a7, tp
                                                  30'd    10647    : data = 32'h    0063DC93    ;    //    srli x25 x7 6      ====        srli s9, t2, 6
                                                  30'd    10648    : data = 32'h    F88E2713    ;    //    slti x14 x28 -120      ====        slti a4, t3, -120
                                                  30'd    10649    : data = 32'h    00E59713    ;    //    slli x14 x11 14      ====        slli a4, a1, 14
                                                  30'd    10650    : data = 32'h    00C9D813    ;    //    srli x16 x19 12      ====        srli a6, s3, 12
                                                  30'd    10651    : data = 32'h    7A45F793    ;    //    andi x15 x11 1956      ====        andi a5, a1, 1956
                                                  30'd    10652    : data = 32'h    01DDF933    ;    //    and x18 x27 x29      ====        and s2, s11, t4
                                                  30'd    10653    : data = 32'h    12540337    ;    //    lui x6 75072      ====        lui t1, 75072
                                                  30'd    10654    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10655    : data = 32'h    016B4833    ;    //    xor x16 x22 x22      ====        xor a6, s6, s6
                                                  30'd    10656    : data = 32'h    C60EB893    ;    //    sltiu x17 x29 -928      ====        sltiu a7, t4, -928
                                                  30'd    10657    : data = 32'h    AD0B7813    ;    //    andi x16 x22 -1328      ====        andi a6, s6, -1328
                                                  30'd    10658    : data = 32'h    416EDD93    ;    //    srai x27 x29 22      ====        srai s11, t4, 22
                                                  30'd    10659    : data = 32'h    4A8CA597    ;    //    auipc x11 305354      ====        auipc a1, 305354
                                                  30'd    10660    : data = 32'h    0193EC33    ;    //    or x24 x7 x25      ====        or s8, t2, s9
                                                  30'd    10661    : data = 32'h    BFD93393    ;    //    sltiu x7 x18 -1027      ====        sltiu t2, s2, -1027
                                                  30'd    10662    : data = 32'h    01EA23B3    ;    //    slt x7 x20 x30      ====        slt t2, s4, t5
                                                  30'd    10663    : data = 32'h    C7948E93    ;    //    addi x29 x9 -903      ====        addi t4, s1, -903
                                                  30'd    10664    : data = 32'h    41D40833    ;    //    sub x16 x8 x29      ====        sub a6, s0, t4
                                                  30'd    10665    : data = 32'h    007F5413    ;    //    srli x8 x30 7      ====        srli s0, t5, 7
                                                  30'd    10666    : data = 32'h    010FF933    ;    //    and x18 x31 x16      ====        and s2, t6, a6
                                                  30'd    10667    : data = 32'h    33035917    ;    //    auipc x18 208949      ====        auipc s2, 208949
                                                  30'd    10668    : data = 32'h    02744313    ;    //    xori x6 x8 39      ====        xori t1, s0, 39
                                                  30'd    10669    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10670    : data = 32'h    408058B3    ;    //    sra x17 x0 x8      ====        sra a7, zero, s0
                                                  30'd    10671    : data = 32'h    00B17BB3    ;    //    and x23 x2 x11      ====        and s7, sp, a1
                                                  30'd    10672    : data = 32'h    00CEA733    ;    //    slt x14 x29 x12      ====        slt a4, t4, a2
                                                  30'd    10673    : data = 32'h    005242B3    ;    //    xor x5 x4 x5      ====        xor t0, tp, t0
                                                  30'd    10674    : data = 32'h    41DA8933    ;    //    sub x18 x21 x29      ====        sub s2, s5, t4
                                                  30'd    10675    : data = 32'h    40FD0FB3    ;    //    sub x31 x26 x15      ====        sub t6, s10, a5
                                                  30'd    10676    : data = 32'h    05147613    ;    //    andi x12 x8 81      ====        andi a2, s0, 81
                                                  30'd    10677    : data = 32'h    00CC41B3    ;    //    xor x3 x24 x12      ====        xor gp, s8, a2
                                                  30'd    10678    : data = 32'h    A4DF8013    ;    //    addi x0 x31 -1459      ====        addi zero, t6, -1459
                                                  30'd    10679    : data = 32'h    00FD1BB3    ;    //    sll x23 x26 x15      ====        sll s7, s10, a5
                                                  30'd    10680    : data = 32'h    418C5A33    ;    //    sra x20 x24 x24      ====        sra s4, s8, s8
                                                  30'd    10681    : data = 32'h    00CF9D13    ;    //    slli x26 x31 12      ====        slli s10, t6, 12
                                                  30'd    10682    : data = 32'h    012D1D13    ;    //    slli x26 x26 18      ====        slli s10, s10, 18
                                                  30'd    10683    : data = 32'h    41205033    ;    //    sra x0 x0 x18      ====        sra zero, zero, s2
                                                  30'd    10684    : data = 32'h    000F8BB3    ;    //    add x23 x31 x0      ====        add s7, t6, zero
                                                  30'd    10685    : data = 32'h    408EDD33    ;    //    sra x26 x29 x8      ====        sra s10, t4, s0
                                                  30'd    10686    : data = 32'h    00EA9693    ;    //    slli x13 x21 14      ====        slli a3, s5, 14
                                                  30'd    10687    : data = 32'h    01044AB3    ;    //    xor x21 x8 x16      ====        xor s5, s0, a6
                                                  30'd    10688    : data = 32'h    018FD193    ;    //    srli x3 x31 24      ====        srli gp, t6, 24
                                                  30'd    10689    : data = 32'h    01E88433    ;    //    add x8 x17 x30      ====        add s0, a7, t5
                                                  30'd    10690    : data = 32'h    E9D6B393    ;    //    sltiu x7 x13 -355      ====        sltiu t2, a3, -355
                                                  30'd    10691    : data = 32'h    45CBD9B7    ;    //    lui x19 285885      ====        lui s3, 285885
                                                  30'd    10692    : data = 32'h    16BB8993    ;    //    addi x19 x23 363      ====        addi s3, s7, 363
                                                  30'd    10693    : data = 32'h    00A1D813    ;    //    srli x16 x3 10      ====        srli a6, gp, 10
                                                  30'd    10694    : data = 32'h    408ADBB3    ;    //    sra x23 x21 x8      ====        sra s7, s5, s0
                                                  30'd    10695    : data = 32'h    412FD013    ;    //    srai x0 x31 18      ====        srai zero, t6, 18
                                                  30'd    10696    : data = 32'h    09D62913    ;    //    slti x18 x12 157      ====        slti s2, a2, 157
                                                  30'd    10697    : data = 32'h    0006AA33    ;    //    slt x20 x13 x0      ====        slt s4, a3, zero
                                                  30'd    10698    : data = 32'h    F2A47B13    ;    //    andi x22 x8 -214      ====        andi s6, s0, -214
                                                  30'd    10699    : data = 32'h    015F1633    ;    //    sll x12 x30 x21      ====        sll a2, t5, s5
                                                  30'd    10700    : data = 32'h    8FB72B13    ;    //    slti x22 x14 -1797      ====        slti s6, a4, -1797
                                                  30'd    10701    : data = 32'h    01E7D493    ;    //    srli x9 x15 30      ====        srli s1, a5, 30
                                                  30'd    10702    : data = 32'h    0081DD13    ;    //    srli x26 x3 8      ====        srli s10, gp, 8
                                                  30'd    10703    : data = 32'h    4119D713    ;    //    srai x14 x19 17      ====        srai a4, s3, 17
                                                  30'd    10704    : data = 32'h    005F20B3    ;    //    slt x1 x30 x5      ====        slt ra, t5, t0
                                                  30'd    10705    : data = 32'h    41E6DDB3    ;    //    sra x27 x13 x30      ====        sra s11, a3, t5
                                                  30'd    10706    : data = 32'h    6F7A7D93    ;    //    andi x27 x20 1783      ====        andi s11, s4, 1783
                                                  30'd    10707    : data = 32'h    414DD333    ;    //    sra x6 x27 x20      ====        sra t1, s11, s4
                                                  30'd    10708    : data = 32'h    0173E733    ;    //    or x14 x7 x23      ====        or a4, t2, s7
                                                  30'd    10709    : data = 32'h    002F39B3    ;    //    sltu x19 x30 x2      ====        sltu s3, t5, sp
                                                  30'd    10710    : data = 32'h    00899093    ;    //    slli x1 x19 8      ====        slli ra, s3, 8
                                                  30'd    10711    : data = 32'h    40B3DD93    ;    //    srai x27 x7 11      ====        srai s11, t2, 11
                                                  30'd    10712    : data = 32'h    409E0333    ;    //    sub x6 x28 x9      ====        sub t1, t3, s1
                                                  30'd    10713    : data = 32'h    0540A713    ;    //    slti x14 x1 84      ====        slti a4, ra, 84
                                                  30'd    10714    : data = 32'h    2F190917    ;    //    auipc x18 192912      ====        auipc s2, 192912
                                                  30'd    10715    : data = 32'h    011ADD33    ;    //    srl x26 x21 x17      ====        srl s10, s5, a7
                                                  30'd    10716    : data = 32'h    CE98C737    ;    //    lui x14 846220      ====        lui a4, 846220
                                                  30'd    10717    : data = 32'h    011136B3    ;    //    sltu x13 x2 x17      ====        sltu a3, sp, a7
                                                  30'd    10718    : data = 32'h    DD262E13    ;    //    slti x28 x12 -558      ====        slti t3, a2, -558
                                                  30'd    10719    : data = 32'h    10184C93    ;    //    xori x25 x16 257      ====        xori s9, a6, 257
                                                  30'd    10720    : data = 32'h    412F82B3    ;    //    sub x5 x31 x18      ====        sub t0, t6, s2
                                                  30'd    10721    : data = 32'h    C815FA97    ;    //    auipc x21 819551      ====        auipc s5, 819551
                                                  30'd    10722    : data = 32'h    0118BD33    ;    //    sltu x26 x17 x17      ====        sltu s10, a7, a7
                                                  30'd    10723    : data = 32'h    EEDF2A13    ;    //    slti x20 x30 -275      ====        slti s4, t5, -275
                                                  30'd    10724    : data = 32'h    01DF4A33    ;    //    xor x20 x30 x29      ====        xor s4, t5, t4
                                                  30'd    10725    : data = 32'h    D33FBD93    ;    //    sltiu x27 x31 -717      ====        sltiu s11, t6, -717
                                                  30'd    10726    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10727    : data = 32'h    00ACF933    ;    //    and x18 x25 x10      ====        and s2, s9, a0
                                                  30'd    10728    : data = 32'h    043F8013    ;    //    addi x0 x31 67      ====        addi zero, t6, 67
                                                  30'd    10729    : data = 32'h    4113DB13    ;    //    srai x22 x7 17      ====        srai s6, t2, 17
                                                  30'd    10730    : data = 32'h    01EDA733    ;    //    slt x14 x27 x30      ====        slt a4, s11, t5
                                                  30'd    10731    : data = 32'h    016318B3    ;    //    sll x17 x6 x22      ====        sll a7, t1, s6
                                                  30'd    10732    : data = 32'h    3C36E113    ;    //    ori x2 x13 963      ====        ori sp, a3, 963
                                                  30'd    10733    : data = 32'h    01D12033    ;    //    slt x0 x2 x29      ====        slt zero, sp, t4
                                                  30'd    10734    : data = 32'h    401A5E13    ;    //    srai x28 x20 1      ====        srai t3, s4, 1
                                                  30'd    10735    : data = 32'h    88CEEE93    ;    //    ori x29 x29 -1908      ====        ori t4, t4, -1908
                                                  30'd    10736    : data = 32'h    00421E33    ;    //    sll x28 x4 x4      ====        sll t3, tp, tp
                                                  30'd    10737    : data = 32'h    01E89D13    ;    //    slli x26 x17 30      ====        slli s10, a7, 30
                                                  30'd    10738    : data = 32'h    0164D413    ;    //    srli x8 x9 22      ====        srli s0, s1, 22
                                                  30'd    10739    : data = 32'h    01AACEB3    ;    //    xor x29 x21 x26      ====        xor t4, s5, s10
                                                  30'd    10740    : data = 32'h    014BFB33    ;    //    and x22 x23 x20      ====        and s6, s7, s4
                                                  30'd    10741    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10742    : data = 32'h    5D81FF93    ;    //    andi x31 x3 1496      ====        andi t6, gp, 1496
                                                  30'd    10743    : data = 32'h    008DE8B3    ;    //    or x17 x27 x8      ====        or a7, s11, s0
                                                  30'd    10744    : data = 32'h    FC343C93    ;    //    sltiu x25 x8 -61      ====        sltiu s9, s0, -61
                                                  30'd    10745    : data = 32'h    006191B3    ;    //    sll x3 x3 x6      ====        sll gp, gp, t1
                                                  30'd    10746    : data = 32'h    001166B3    ;    //    or x13 x2 x1      ====        or a3, sp, ra
                                                  30'd    10747    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10748    : data = 32'h    89A27597    ;    //    auipc x11 563751      ====        auipc a1, 563751
                                                  30'd    10749    : data = 32'h    F9310917    ;    //    auipc x18 1020688      ====        auipc s2, 1020688
                                                  30'd    10750    : data = 32'h    0050CC33    ;    //    xor x24 x1 x5      ====        xor s8, ra, t0
                                                  30'd    10751    : data = 32'h    00D879B3    ;    //    and x19 x16 x13      ====        and s3, a6, a3
                                                  30'd    10752    : data = 32'h    CBF70F93    ;    //    addi x31 x14 -833      ====        addi t6, a4, -833
                                                  30'd    10753    : data = 32'h    F7BCDF97    ;    //    auipc x31 1014733      ====        auipc t6, 1014733
                                                  30'd    10754    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10755    : data = 32'h    40558BB3    ;    //    sub x23 x11 x5      ====        sub s7, a1, t0
                                                  30'd    10756    : data = 32'h    2A64A797    ;    //    auipc x15 173642      ====        auipc a5, 173642
                                                  30'd    10757    : data = 32'h    01488CB3    ;    //    add x25 x17 x20      ====        add s9, a7, s4
                                                  30'd    10758    : data = 32'h    40375B33    ;    //    sra x22 x14 x3      ====        sra s6, a4, gp
                                                  30'd    10759    : data = 32'h    009677B3    ;    //    and x15 x12 x9      ====        and a5, a2, s1
                                                  30'd    10760    : data = 32'h    B1F93593    ;    //    sltiu x11 x18 -1249      ====        sltiu a1, s2, -1249
                                                  30'd    10761    : data = 32'h    2B03B693    ;    //    sltiu x13 x7 688      ====        sltiu a3, t2, 688
                                                  30'd    10762    : data = 32'h    E0423693    ;    //    sltiu x13 x4 -508      ====        sltiu a3, tp, -508
                                                  30'd    10763    : data = 32'h    D8900B93    ;    //    addi x23 x0 -631      ====        addi s7, zero, -631
                                                  30'd    10764    : data = 32'h    015AA8B3    ;    //    slt x17 x21 x21      ====        slt a7, s5, s5
                                                  30'd    10765    : data = 32'h    0110C1B3    ;    //    xor x3 x1 x17      ====        xor gp, ra, a7
                                                  30'd    10766    : data = 32'h    006D59B3    ;    //    srl x19 x26 x6      ====        srl s3, s10, t1
                                                  30'd    10767    : data = 32'h    01E26433    ;    //    or x8 x4 x30      ====        or s0, tp, t5
                                                  30'd    10768    : data = 32'h    50264493    ;    //    xori x9 x12 1282      ====        xori s1, a2, 1282
                                                  30'd    10769    : data = 32'h    00EDCB33    ;    //    xor x22 x27 x14      ====        xor s6, s11, a4
                                                  30'd    10770    : data = 32'h    F8564493    ;    //    xori x9 x12 -123      ====        xori s1, a2, -123
                                                  30'd    10771    : data = 32'h    423964B7    ;    //    lui x9 271254      ====        lui s1, 271254
                                                  30'd    10772    : data = 32'h    00BF7EB3    ;    //    and x29 x30 x11      ====        and t4, t5, a1
                                                  30'd    10773    : data = 32'h    01AD02B3    ;    //    add x5 x26 x26      ====        add t0, s10, s10
                                                  30'd    10774    : data = 32'h    01709413    ;    //    slli x8 x1 23      ====        slli s0, ra, 23
                                                  30'd    10775    : data = 32'h    00AFC6B3    ;    //    xor x13 x31 x10      ====        xor a3, t6, a0
                                                  30'd    10776    : data = 32'h    41B0D713    ;    //    srai x14 x1 27      ====        srai a4, ra, 27
                                                  30'd    10777    : data = 32'h    85EAD937    ;    //    lui x18 548525      ====        lui s2, 548525
                                                  30'd    10778    : data = 32'h    015705B3    ;    //    add x11 x14 x21      ====        add a1, a4, s5
                                                  30'd    10779    : data = 32'h    EC4B4193    ;    //    xori x3 x22 -316      ====        xori gp, s6, -316
                                                  30'd    10780    : data = 32'h    00251CB3    ;    //    sll x25 x10 x2      ====        sll s9, a0, sp
                                                  30'd    10781    : data = 32'h    40095613    ;    //    srai x12 x18 0      ====        srai a2, s2, 0
                                                  30'd    10782    : data = 32'h    00809D13    ;    //    slli x26 x1 8      ====        slli s10, ra, 8
                                                  30'd    10783    : data = 32'h    BEF69737    ;    //    lui x14 782185      ====        lui a4, 782185
                                                  30'd    10784    : data = 32'h    7D0D2D13    ;    //    slti x26 x26 2000      ====        slti s10, s10, 2000
                                                  30'd    10785    : data = 32'h    0E97EE97    ;    //    auipc x29 59774      ====        auipc t4, 59774
                                                  30'd    10786    : data = 32'h    4EADE293    ;    //    ori x5 x27 1258      ====        ori t0, s11, 1258
                                                  30'd    10787    : data = 32'h    A313A417    ;    //    auipc x8 667962      ====        auipc s0, 667962
                                                  30'd    10788    : data = 32'h    011A5F93    ;    //    srli x31 x20 17      ====        srli t6, s4, 17
                                                  30'd    10789    : data = 32'h    416ADB33    ;    //    sra x22 x21 x22      ====        sra s6, s5, s6
                                                  30'd    10790    : data = 32'h    01AE1133    ;    //    sll x2 x28 x26      ====        sll sp, t3, s10
                                                  30'd    10791    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10792    : data = 32'h    00928733    ;    //    add x14 x5 x9      ====        add a4, t0, s1
                                                  30'd    10793    : data = 32'h    00321113    ;    //    slli x2 x4 3      ====        slli sp, tp, 3
                                                  30'd    10794    : data = 32'h    013A9733    ;    //    sll x14 x21 x19      ====        sll a4, s5, s3
                                                  30'd    10795    : data = 32'h    91AD2313    ;    //    slti x6 x26 -1766      ====        slti t1, s10, -1766
                                                  30'd    10796    : data = 32'h    86A70B93    ;    //    addi x23 x14 -1942      ====        addi s7, a4, -1942
                                                  30'd    10797    : data = 32'h    0012FD33    ;    //    and x26 x5 x1      ====        and s10, t0, ra
                                                  30'd    10798    : data = 32'h    00CA2EB3    ;    //    slt x29 x20 x12      ====        slt t4, s4, a2
                                                  30'd    10799    : data = 32'h    40680733    ;    //    sub x14 x16 x6      ====        sub a4, a6, t1
                                                  30'd    10800    : data = 32'h    0085BCB3    ;    //    sltu x25 x11 x8      ====        sltu s9, a1, s0
                                                  30'd    10801    : data = 32'h    016E3DB3    ;    //    sltu x27 x28 x22      ====        sltu s11, t3, s6
                                                  30'd    10802    : data = 32'h    40425413    ;    //    srai x8 x4 4      ====        srai s0, tp, 4
                                                  30'd    10803    : data = 32'h    621CDC17    ;    //    auipc x24 401869      ====        auipc s8, 401869
                                                  30'd    10804    : data = 32'h    7741A393    ;    //    slti x7 x3 1908      ====        slti t2, gp, 1908
                                                  30'd    10805    : data = 32'h    01815313    ;    //    srli x6 x2 24      ====        srli t1, sp, 24
                                                  30'd    10806    : data = 32'h    4145D9B3    ;    //    sra x19 x11 x20      ====        sra s3, a1, s4
                                                  30'd    10807    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10808    : data = 32'h    00A0DEB3    ;    //    srl x29 x1 x10      ====        srl t4, ra, a0
                                                  30'd    10809    : data = 32'h    01CEB9B3    ;    //    sltu x19 x29 x28      ====        sltu s3, t4, t3
                                                  30'd    10810    : data = 32'h    00B71733    ;    //    sll x14 x14 x11      ====        sll a4, a4, a1
                                                  30'd    10811    : data = 32'h    00B4E933    ;    //    or x18 x9 x11      ====        or s2, s1, a1
                                                  30'd    10812    : data = 32'h    CD8CB413    ;    //    sltiu x8 x25 -808      ====        sltiu s0, s9, -808
                                                  30'd    10813    : data = 32'h    00E0CE33    ;    //    xor x28 x1 x14      ====        xor t3, ra, a4
                                                  30'd    10814    : data = 32'h    0106D093    ;    //    srli x1 x13 16      ====        srli ra, a3, 16
                                                  30'd    10815    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10816    : data = 32'h    A014AA93    ;    //    slti x21 x9 -1535      ====        slti s5, s1, -1535
                                                  30'd    10817    : data = 32'h    F8D683B7    ;    //    lui x7 1019240      ====        lui t2, 1019240
                                                  30'd    10818    : data = 32'h    00180133    ;    //    add x2 x16 x1      ====        add sp, a6, ra
                                                  30'd    10819    : data = 32'h    4060D0B3    ;    //    sra x1 x1 x6      ====        sra ra, ra, t1
                                                  30'd    10820    : data = 32'h    2F4E2B93    ;    //    slti x23 x28 756      ====        slti s7, t3, 756
                                                  30'd    10821    : data = 32'h    00245813    ;    //    srli x16 x8 2      ====        srli a6, s0, 2
                                                  30'd    10822    : data = 32'h    40B95113    ;    //    srai x2 x18 11      ====        srai sp, s2, 11
                                                  30'd    10823    : data = 32'h    416A53B3    ;    //    sra x7 x20 x22      ====        sra t2, s4, s6
                                                  30'd    10824    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10825    : data = 32'h    F5EFAD93    ;    //    slti x27 x31 -162      ====        slti s11, t6, -162
                                                  30'd    10826    : data = 32'h    014D2E33    ;    //    slt x28 x26 x20      ====        slt t3, s10, s4
                                                  30'd    10827    : data = 32'h    4D98B113    ;    //    sltiu x2 x17 1241      ====        sltiu sp, a7, 1241
                                                  30'd    10828    : data = 32'h    0048D7B3    ;    //    srl x15 x17 x4      ====        srl a5, a7, tp
                                                  30'd    10829    : data = 32'h    41465633    ;    //    sra x12 x12 x20      ====        sra a2, a2, s4
                                                  30'd    10830    : data = 32'h    52DCE293    ;    //    ori x5 x25 1325      ====        ori t0, s9, 1325
                                                  30'd    10831    : data = 32'h    01065F93    ;    //    srli x31 x12 16      ====        srli t6, a2, 16
                                                  30'd    10832    : data = 32'h    015AA4B3    ;    //    slt x9 x21 x21      ====        slt s1, s5, s5
                                                  30'd    10833    : data = 32'h    1D8F6693    ;    //    ori x13 x30 472      ====        ori a3, t5, 472
                                                  30'd    10834    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10835    : data = 32'h    61A07E93    ;    //    andi x29 x0 1562      ====        andi t4, zero, 1562
                                                  30'd    10836    : data = 32'h    41FBD293    ;    //    srai x5 x23 31      ====        srai t0, s7, 31
                                                  30'd    10837    : data = 32'h    00065093    ;    //    srli x1 x12 0      ====        srli ra, a2, 0
                                                  30'd    10838    : data = 32'h    AD286113    ;    //    ori x2 x16 -1326      ====        ori sp, a6, -1326
                                                  30'd    10839    : data = 32'h    00FA41B3    ;    //    xor x3 x20 x15      ====        xor gp, s4, a5
                                                  30'd    10840    : data = 32'h    8062E613    ;    //    ori x12 x5 -2042      ====        ori a2, t0, -2042
                                                  30'd    10841    : data = 32'h    9EE34613    ;    //    xori x12 x6 -1554      ====        xori a2, t1, -1554
                                                  30'd    10842    : data = 32'h    01061693    ;    //    slli x13 x12 16      ====        slli a3, a2, 16
                                                  30'd    10843    : data = 32'h    019A61B3    ;    //    or x3 x20 x25      ====        or gp, s4, s9
                                                  30'd    10844    : data = 32'h    AD2A0593    ;    //    addi x11 x20 -1326      ====        addi a1, s4, -1326
                                                  30'd    10845    : data = 32'h    419E8BB3    ;    //    sub x23 x29 x25      ====        sub s7, t4, s9
                                                  30'd    10846    : data = 32'h    0122E633    ;    //    or x12 x5 x18      ====        or a2, t0, s2
                                                  30'd    10847    : data = 32'h    00899FB3    ;    //    sll x31 x19 x8      ====        sll t6, s3, s0
                                                  30'd    10848    : data = 32'h    413A5633    ;    //    sra x12 x20 x19      ====        sra a2, s4, s3
                                                  30'd    10849    : data = 32'h    F9DA6837    ;    //    lui x16 1023398      ====        lui a6, 1023398
                                                  30'd    10850    : data = 32'h    004E9A13    ;    //    slli x20 x29 4      ====        slli s4, t4, 4
                                                  30'd    10851    : data = 32'h    D163F713    ;    //    andi x14 x7 -746      ====        andi a4, t2, -746
                                                  30'd    10852    : data = 32'h    47504F93    ;    //    xori x31 x0 1141      ====        xori t6, zero, 1141
                                                  30'd    10853    : data = 32'h    00B8A0B3    ;    //    slt x1 x17 x11      ====        slt ra, a7, a1
                                                  30'd    10854    : data = 32'h    00438133    ;    //    add x2 x7 x4      ====        add sp, t2, tp
                                                  30'd    10855    : data = 32'h    01D55E33    ;    //    srl x28 x10 x29      ====        srl t3, a0, t4
                                                  30'd    10856    : data = 32'h    01F55613    ;    //    srli x12 x10 31      ====        srli a2, a0, 31
                                                  30'd    10857    : data = 32'h    010C95B3    ;    //    sll x11 x25 x16      ====        sll a1, s9, a6
                                                  30'd    10858    : data = 32'h    00A728B3    ;    //    slt x17 x14 x10      ====        slt a7, a4, a0
                                                  30'd    10859    : data = 32'h    006837B3    ;    //    sltu x15 x16 x6      ====        sltu a5, a6, t1
                                                  30'd    10860    : data = 32'h    35EFB0B7    ;    //    lui x1 220923      ====        lui ra, 220923
                                                  30'd    10861    : data = 32'h    01A5DC13    ;    //    srli x24 x11 26      ====        srli s8, a1, 26
                                                  30'd    10862    : data = 32'h    DDBDD797    ;    //    auipc x15 908253      ====        auipc a5, 908253
                                                  30'd    10863    : data = 32'h    32C19A37    ;    //    lui x20 207897      ====        lui s4, 207897
                                                  30'd    10864    : data = 32'h    014D39B3    ;    //    sltu x19 x26 x20      ====        sltu s3, s10, s4
                                                  30'd    10865    : data = 32'h    00A90033    ;    //    add x0 x18 x10      ====        add zero, s2, a0
                                                  30'd    10866    : data = 32'h    57297D13    ;    //    andi x26 x18 1394      ====        andi s10, s2, 1394
                                                  30'd    10867    : data = 32'h    E5A9BB93    ;    //    sltiu x23 x19 -422      ====        sltiu s7, s3, -422
                                                  30'd    10868    : data = 32'h    01A2B2B3    ;    //    sltu x5 x5 x26      ====        sltu t0, t0, s10
                                                  30'd    10869    : data = 32'h    18C30113    ;    //    addi x2 x6 396      ====        addi sp, t1, 396
                                                  30'd    10870    : data = 32'h    01AB66B3    ;    //    or x13 x22 x26      ====        or a3, s6, s10
                                                  30'd    10871    : data = 32'h    B73AE693    ;    //    ori x13 x21 -1165      ====        ori a3, s5, -1165
                                                  30'd    10872    : data = 32'h    4105D613    ;    //    srai x12 x11 16      ====        srai a2, a1, 16
                                                  30'd    10873    : data = 32'h    01773CB3    ;    //    sltu x25 x14 x23      ====        sltu s9, a4, s7
                                                  30'd    10874    : data = 32'h    00A6ECB3    ;    //    or x25 x13 x10      ====        or s9, a3, a0
                                                  30'd    10875    : data = 32'h    BA4F37B7    ;    //    lui x15 763123      ====        lui a5, 763123
                                                  30'd    10876    : data = 32'h    0074B3B3    ;    //    sltu x7 x9 x7      ====        sltu t2, s1, t2
                                                  30'd    10877    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10878    : data = 32'h    00CF7433    ;    //    and x8 x30 x12      ====        and s0, t5, a2
                                                  30'd    10879    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10880    : data = 32'h    83B4FD93    ;    //    andi x27 x9 -1989      ====        andi s11, s1, -1989
                                                  30'd    10881    : data = 32'h    FE2B0D93    ;    //    addi x27 x22 -30      ====        addi s11, s6, -30
                                                  30'd    10882    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10883    : data = 32'h    00D841B3    ;    //    xor x3 x16 x13      ====        xor gp, a6, a3
                                                  30'd    10884    : data = 32'h    010C8D33    ;    //    add x26 x25 x16      ====        add s10, s9, a6
                                                  30'd    10885    : data = 32'h    40465033    ;    //    sra x0 x12 x4      ====        sra zero, a2, tp
                                                  30'd    10886    : data = 32'h    1B790613    ;    //    addi x12 x18 439      ====        addi a2, s2, 439
                                                  30'd    10887    : data = 32'h    40CA0E33    ;    //    sub x28 x20 x12      ====        sub t3, s4, a2
                                                  30'd    10888    : data = 32'h    008B9933    ;    //    sll x18 x23 x8      ====        sll s2, s7, s0
                                                  30'd    10889    : data = 32'h    011C03B3    ;    //    add x7 x24 x17      ====        add t2, s8, a7
                                                  30'd    10890    : data = 32'h    40C4D5B3    ;    //    sra x11 x9 x12      ====        sra a1, s1, a2
                                                  30'd    10891    : data = 32'h    00C2C733    ;    //    xor x14 x5 x12      ====        xor a4, t0, a2
                                                  30'd    10892    : data = 32'h    01F61D13    ;    //    slli x26 x12 31      ====        slli s10, a2, 31
                                                  30'd    10893    : data = 32'h    005CBC33    ;    //    sltu x24 x25 x5      ====        sltu s8, s9, t0
                                                  30'd    10894    : data = 32'h    37A42E13    ;    //    slti x28 x8 890      ====        slti t3, s0, 890
                                                  30'd    10895    : data = 32'h    13769597    ;    //    auipc x11 79721      ====        auipc a1, 79721
                                                  30'd    10896    : data = 32'h    009889B3    ;    //    add x19 x17 x9      ====        add s3, a7, s1
                                                  30'd    10897    : data = 32'h    8795B397    ;    //    auipc x7 555355      ====        auipc t2, 555355
                                                  30'd    10898    : data = 32'h    623E8B13    ;    //    addi x22 x29 1571      ====        addi s6, t4, 1571
                                                  30'd    10899    : data = 32'h    01A3DA33    ;    //    srl x20 x7 x26      ====        srl s4, t2, s10
                                                  30'd    10900    : data = 32'h    015960B3    ;    //    or x1 x18 x21      ====        or ra, s2, s5
                                                  30'd    10901    : data = 32'h    405AD933    ;    //    sra x18 x21 x5      ====        sra s2, s5, t0
                                                  30'd    10902    : data = 32'h    9C6D0893    ;    //    addi x17 x26 -1594      ====        addi a7, s10, -1594
                                                  30'd    10903    : data = 32'h    0018CEB3    ;    //    xor x29 x17 x1      ====        xor t4, a7, ra
                                                  30'd    10904    : data = 32'h    7AE5AB13    ;    //    slti x22 x11 1966      ====        slti s6, a1, 1966
                                                  30'd    10905    : data = 32'h    72424413    ;    //    xori x8 x4 1828      ====        xori s0, tp, 1828
                                                  30'd    10906    : data = 32'h    00B10033    ;    //    add x0 x2 x11      ====        add zero, sp, a1
                                                  30'd    10907    : data = 32'h    F6D08D93    ;    //    addi x27 x1 -147      ====        addi s11, ra, -147
                                                  30'd    10908    : data = 32'h    009AC833    ;    //    xor x16 x21 x9      ====        xor a6, s5, s1
                                                  30'd    10909    : data = 32'h    006FC1B3    ;    //    xor x3 x31 x6      ====        xor gp, t6, t1
                                                  30'd    10910    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10911    : data = 32'h    41F95813    ;    //    srai x16 x18 31      ====        srai a6, s2, 31
                                                  30'd    10912    : data = 32'h    B6256D13    ;    //    ori x26 x10 -1182      ====        ori s10, a0, -1182
                                                  30'd    10913    : data = 32'h    019A6C33    ;    //    or x24 x20 x25      ====        or s8, s4, s9
                                                  30'd    10914    : data = 32'h    013BB033    ;    //    sltu x0 x23 x19      ====        sltu zero, s7, s3
                                                  30'd    10915    : data = 32'h    41BFD033    ;    //    sra x0 x31 x27      ====        sra zero, t6, s11
                                                  30'd    10916    : data = 32'h    DDEA6B93    ;    //    ori x23 x20 -546      ====        ori s7, s4, -546
                                                  30'd    10917    : data = 32'h    2B18EA13    ;    //    ori x20 x17 689      ====        ori s4, a7, 689
                                                  30'd    10918    : data = 32'h    00B66E33    ;    //    or x28 x12 x11      ====        or t3, a2, a1
                                                  30'd    10919    : data = 32'h    416AD393    ;    //    srai x7 x21 22      ====        srai t2, s5, 22
                                                  30'd    10920    : data = 32'h    01908BB3    ;    //    add x23 x1 x25      ====        add s7, ra, s9
                                                  30'd    10921    : data = 32'h    74CECA93    ;    //    xori x21 x29 1868      ====        xori s5, t4, 1868
                                                  30'd    10922    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10923    : data = 32'h    798E3193    ;    //    sltiu x3 x28 1944      ====        sltiu gp, t3, 1944
                                                  30'd    10924    : data = 32'h    40C68433    ;    //    sub x8 x13 x12      ====        sub s0, a3, a2
                                                  30'd    10925    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10926    : data = 32'h    0097C2B3    ;    //    xor x5 x15 x9      ====        xor t0, a5, s1
                                                  30'd    10927    : data = 32'h    00F5F1B3    ;    //    and x3 x11 x15      ====        and gp, a1, a5
                                                  30'd    10928    : data = 32'h    B1F26E13    ;    //    ori x28 x4 -1249      ====        ori t3, tp, -1249
                                                  30'd    10929    : data = 32'h    4148DE13    ;    //    srai x28 x17 20      ====        srai t3, a7, 20
                                                  30'd    10930    : data = 32'h    41870FB3    ;    //    sub x31 x14 x24      ====        sub t6, a4, s8
                                                  30'd    10931    : data = 32'h    EFF54A93    ;    //    xori x21 x10 -257      ====        xori s5, a0, -257
                                                  30'd    10932    : data = 32'h    001C1C93    ;    //    slli x25 x24 1      ====        slli s9, s8, 1
                                                  30'd    10933    : data = 32'h    D8439B37    ;    //    lui x22 885817      ====        lui s6, 885817
                                                  30'd    10934    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10935    : data = 32'h    00541D33    ;    //    sll x26 x8 x5      ====        sll s10, s0, t0
                                                  30'd    10936    : data = 32'h    40F4D633    ;    //    sra x12 x9 x15      ====        sra a2, s1, a5
                                                  30'd    10937    : data = 32'h    BC086D17    ;    //    auipc x26 770182      ====        auipc s10, 770182
                                                  30'd    10938    : data = 32'h    003E4E33    ;    //    xor x28 x28 x3      ====        xor t3, t3, gp
                                                  30'd    10939    : data = 32'h    01DD9D33    ;    //    sll x26 x27 x29      ====        sll s10, s11, t4
                                                  30'd    10940    : data = 32'h    00F39133    ;    //    sll x2 x7 x15      ====        sll sp, t2, a5
                                                  30'd    10941    : data = 32'h    9B1E7413    ;    //    andi x8 x28 -1615      ====        andi s0, t3, -1615
                                                  30'd    10942    : data = 32'h    40BFDB93    ;    //    srai x23 x31 11      ====        srai s7, t6, 11
                                                  30'd    10943    : data = 32'h    401CD413    ;    //    srai x8 x25 1      ====        srai s0, s9, 1
                                                  30'd    10944    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10945    : data = 32'h    418D8633    ;    //    sub x12 x27 x24      ====        sub a2, s11, s8
                                                  30'd    10946    : data = 32'h    401B8BB3    ;    //    sub x23 x23 x1      ====        sub s7, s7, ra
                                                  30'd    10947    : data = 32'h    010B7D33    ;    //    and x26 x22 x16      ====        and s10, s6, a6
                                                  30'd    10948    : data = 32'h    40F10B33    ;    //    sub x22 x2 x15      ====        sub s6, sp, a5
                                                  30'd    10949    : data = 32'h    00E83BB3    ;    //    sltu x23 x16 x14      ====        sltu s7, a6, a4
                                                  30'd    10950    : data = 32'h    5F008A93    ;    //    addi x21 x1 1520      ====        addi s5, ra, 1520
                                                  30'd    10951    : data = 32'h    41885493    ;    //    srai x9 x16 24      ====        srai s1, a6, 24
                                                  30'd    10952    : data = 32'h    00E8F133    ;    //    and x2 x17 x14      ====        and sp, a7, a4
                                                  30'd    10953    : data = 32'h    00F0D413    ;    //    srli x8 x1 15      ====        srli s0, ra, 15
                                                  30'd    10954    : data = 32'h    9AE7B193    ;    //    sltiu x3 x15 -1618      ====        sltiu gp, a5, -1618
                                                  30'd    10955    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10956    : data = 32'h    17AC6D17    ;    //    auipc x26 96966      ====        auipc s10, 96966
                                                  30'd    10957    : data = 32'h    014C9693    ;    //    slli x13 x25 20      ====        slli a3, s9, 20
                                                  30'd    10958    : data = 32'h    40ED5E13    ;    //    srai x28 x26 14      ====        srai t3, s10, 14
                                                  30'd    10959    : data = 32'h    8FFCF193    ;    //    andi x3 x25 -1793      ====        andi gp, s9, -1793
                                                  30'd    10960    : data = 32'h    41128B33    ;    //    sub x22 x5 x17      ====        sub s6, t0, a7
                                                  30'd    10961    : data = 32'h    5DFD2993    ;    //    slti x19 x26 1503      ====        slti s3, s10, 1503
                                                  30'd    10962    : data = 32'h    011A67B3    ;    //    or x15 x20 x17      ====        or a5, s4, a7
                                                  30'd    10963    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10964    : data = 32'h    98440B13    ;    //    addi x22 x8 -1660      ====        addi s6, s0, -1660
                                                  30'd    10965    : data = 32'h    07C61EB7    ;    //    lui x29 31841      ====        lui t4, 31841
                                                  30'd    10966    : data = 32'h    40D102B3    ;    //    sub x5 x2 x13      ====        sub t0, sp, a3
                                                  30'd    10967    : data = 32'h    00BA9B33    ;    //    sll x22 x21 x11      ====        sll s6, s5, a1
                                                  30'd    10968    : data = 32'h    0096DD33    ;    //    srl x26 x13 x9      ====        srl s10, a3, s1
                                                  30'd    10969    : data = 32'h    00E3F733    ;    //    and x14 x7 x14      ====        and a4, t2, a4
                                                  30'd    10970    : data = 32'h    00BB4633    ;    //    xor x12 x22 x11      ====        xor a2, s6, a1
                                                  30'd    10971    : data = 32'h    00FCAD33    ;    //    slt x26 x25 x15      ====        slt s10, s9, a5
                                                  30'd    10972    : data = 32'h    D15B6113    ;    //    ori x2 x22 -747      ====        ori sp, s6, -747
                                                  30'd    10973    : data = 32'h    01A83D33    ;    //    sltu x26 x16 x26      ====        sltu s10, a6, s10
                                                  30'd    10974    : data = 32'h    401E8933    ;    //    sub x18 x29 x1      ====        sub s2, t4, ra
                                                  30'd    10975    : data = 32'h    01552933    ;    //    slt x18 x10 x21      ====        slt s2, a0, s5
                                                  30'd    10976    : data = 32'h    01A6C733    ;    //    xor x14 x13 x26      ====        xor a4, a3, s10
                                                  30'd    10977    : data = 32'h    59F4A413    ;    //    slti x8 x9 1439      ====        slti s0, s1, 1439
                                                  30'd    10978    : data = 32'h    01D5D293    ;    //    srli x5 x11 29      ====        srli t0, a1, 29
                                                  30'd    10979    : data = 32'h    01A08D33    ;    //    add x26 x1 x26      ====        add s10, ra, s10
                                                  30'd    10980    : data = 32'h    00C58633    ;    //    add x12 x11 x12      ====        add a2, a1, a2
                                                  30'd    10981    : data = 32'h    78A8CD93    ;    //    xori x27 x17 1930      ====        xori s11, a7, 1930
                                                  30'd    10982    : data = 32'h    66BD3C17    ;    //    auipc x24 420819      ====        auipc s8, 420819
                                                  30'd    10983    : data = 32'h    A8F8DA17    ;    //    auipc x20 692109      ====        auipc s4, 692109
                                                  30'd    10984    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    10985    : data = 32'h    00E39013    ;    //    slli x0 x7 14      ====        slli zero, t2, 14
                                                  30'd    10986    : data = 32'h    0141BEB3    ;    //    sltu x29 x3 x20      ====        sltu t4, gp, s4
                                                  30'd    10987    : data = 32'h    01C7E133    ;    //    or x2 x15 x28      ====        or sp, a5, t3
                                                  30'd    10988    : data = 32'h    C1363093    ;    //    sltiu x1 x12 -1005      ====        sltiu ra, a2, -1005
                                                  30'd    10989    : data = 32'h    828A7313    ;    //    andi x6 x20 -2008      ====        andi t1, s4, -2008
                                                  30'd    10990    : data = 32'h    4047DD13    ;    //    srai x26 x15 4      ====        srai s10, a5, 4
                                                  30'd    10991    : data = 32'h    62762B97    ;    //    auipc x23 403298      ====        auipc s7, 403298
                                                  30'd    10992    : data = 32'h    01D89B93    ;    //    slli x23 x17 29      ====        slli s7, a7, 29
                                                  30'd    10993    : data = 32'h    01A58AB3    ;    //    add x21 x11 x26      ====        add s5, a1, s10
                                                  30'd    10994    : data = 32'h    00E2B733    ;    //    sltu x14 x5 x14      ====        sltu a4, t0, a4
                                                  30'd    10995    : data = 32'h    53DA0997    ;    //    auipc x19 343456      ====        auipc s3, 343456
                                                  30'd    10996    : data = 32'h    C67F7D13    ;    //    andi x26 x30 -921      ====        andi s10, t5, -921
                                                  30'd    10997    : data = 32'h    79258993    ;    //    addi x19 x11 1938      ====        addi s3, a1, 1938
                                                  30'd    10998    : data = 32'h    3A707193    ;    //    andi x3 x0 935      ====        andi gp, zero, 935
                                                  30'd    10999    : data = 32'h    01847933    ;    //    and x18 x8 x24      ====        and s2, s0, s8
                                                  30'd    11000    : data = 32'h    01B7ABB3    ;    //    slt x23 x15 x27      ====        slt s7, a5, s11
                                                  30'd    11001    : data = 32'h    0012D013    ;    //    srli x0 x5 1      ====        srli zero, t0, 1
                                                  30'd    11002    : data = 32'h    005EB5B3    ;    //    sltu x11 x29 x5      ====        sltu a1, t4, t0
                                                  30'd    11003    : data = 32'h    00C11733    ;    //    sll x14 x2 x12      ====        sll a4, sp, a2
                                                  30'd    11004    : data = 32'h    8900AE13    ;    //    slti x28 x1 -1904      ====        slti t3, ra, -1904
                                                  30'd    11005    : data = 32'h    CB402713    ;    //    slti x14 x0 -844      ====        slti a4, zero, -844
                                                  30'd    11006    : data = 32'h    019713B3    ;    //    sll x7 x14 x25      ====        sll t2, a4, s9
                                                  30'd    11007    : data = 32'h    01C20EB3    ;    //    add x29 x4 x28      ====        add t4, tp, t3
                                                  30'd    11008    : data = 32'h    01E41933    ;    //    sll x18 x8 x30      ====        sll s2, s0, t5
                                                  30'd    11009    : data = 32'h    009D1FB3    ;    //    sll x31 x26 x9      ====        sll t6, s10, s1
                                                  30'd    11010    : data = 32'h    0192E5B3    ;    //    or x11 x5 x25      ====        or a1, t0, s9
                                                  30'd    11011    : data = 32'h    012A5D13    ;    //    srli x26 x20 18      ====        srli s10, s4, 18
                                                  30'd    11012    : data = 32'h    00561C13    ;    //    slli x24 x12 5      ====        slli s8, a2, 5
                                                  30'd    11013    : data = 32'h    00DA3D33    ;    //    sltu x26 x20 x13      ====        sltu s10, s4, a3
                                                  30'd    11014    : data = 32'h    00A15713    ;    //    srli x14 x2 10      ====        srli a4, sp, 10
                                                  30'd    11015    : data = 32'h    6A1D7C13    ;    //    andi x24 x26 1697      ====        andi s8, s10, 1697
                                                  30'd    11016    : data = 32'h    40EED433    ;    //    sra x8 x29 x14      ====        sra s0, t4, a4
                                                  30'd    11017    : data = 32'h    01333633    ;    //    sltu x12 x6 x19      ====        sltu a2, t1, s3
                                                  30'd    11018    : data = 32'h    06D63B13    ;    //    sltiu x22 x12 109      ====        sltiu s6, a2, 109
                                                  30'd    11019    : data = 32'h    A5CF3913    ;    //    sltiu x18 x30 -1444      ====        sltiu s2, t5, -1444
                                                  30'd    11020    : data = 32'h    01891813    ;    //    slli x16 x18 24      ====        slli a6, s2, 24
                                                  30'd    11021    : data = 32'h    F43B7BB7    ;    //    lui x23 1000375      ====        lui s7, 1000375
                                                  30'd    11022    : data = 32'h    00100CB3    ;    //    add x25 x0 x1      ====        add s9, zero, ra
                                                  30'd    11023    : data = 32'h    0180ED33    ;    //    or x26 x1 x24      ====        or s10, ra, s8
                                                  30'd    11024    : data = 32'h    012F1C93    ;    //    slli x25 x30 18      ====        slli s9, t5, 18
                                                  30'd    11025    : data = 32'h    01D12733    ;    //    slt x14 x2 x29      ====        slt a4, sp, t4
                                                  30'd    11026    : data = 32'h    012FB2B3    ;    //    sltu x5 x31 x18      ====        sltu t0, t6, s2
                                                  30'd    11027    : data = 32'h    6B81B293    ;    //    sltiu x5 x3 1720      ====        sltiu t0, gp, 1720
                                                  30'd    11028    : data = 32'h    0205E013    ;    //    ori x0 x11 32      ====        ori zero, a1, 32
                                                  30'd    11029    : data = 32'h    00441B93    ;    //    slli x23 x8 4      ====        slli s7, s0, 4
                                                  30'd    11030    : data = 32'h    6C2D3413    ;    //    sltiu x8 x26 1730      ====        sltiu s0, s10, 1730
                                                  30'd    11031    : data = 32'h    014917B3    ;    //    sll x15 x18 x20      ====        sll a5, s2, s4
                                                  30'd    11032    : data = 32'h    00A91693    ;    //    slli x13 x18 10      ====        slli a3, s2, 10
                                                  30'd    11033    : data = 32'h    0040E333    ;    //    or x6 x1 x4      ====        or t1, ra, tp
                                                  30'd    11034    : data = 32'h    54217E93    ;    //    andi x29 x2 1346      ====        andi t4, sp, 1346
                                                  30'd    11035    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11036    : data = 32'h    5B5604B7    ;    //    lui x9 374112      ====        lui s1, 374112
                                                  30'd    11037    : data = 32'h    634D0313    ;    //    addi x6 x26 1588      ====        addi t1, s10, 1588
                                                  30'd    11038    : data = 32'h    50904013    ;    //    xori x0 x0 1289      ====        xori zero, zero, 1289
                                                  30'd    11039    : data = 32'h    00A136B3    ;    //    sltu x13 x2 x10      ====        sltu a3, sp, a0
                                                  30'd    11040    : data = 32'h    00FC2A33    ;    //    slt x20 x24 x15      ====        slt s4, s8, a5
                                                  30'd    11041    : data = 32'h    74756D93    ;    //    ori x27 x10 1863      ====        ori s11, a0, 1863
                                                  30'd    11042    : data = 32'h    C0C74C93    ;    //    xori x25 x14 -1012      ====        xori s9, a4, -1012
                                                  30'd    11043    : data = 32'h    41E45833    ;    //    sra x16 x8 x30      ====        sra a6, s0, t5
                                                  30'd    11044    : data = 32'h    0123A9B3    ;    //    slt x19 x7 x18      ====        slt s3, t2, s2
                                                  30'd    11045    : data = 32'h    01771113    ;    //    slli x2 x14 23      ====        slli sp, a4, 23
                                                  30'd    11046    : data = 32'h    0118D013    ;    //    srli x0 x17 17      ====        srli zero, a7, 17
                                                  30'd    11047    : data = 32'h    01E2E433    ;    //    or x8 x5 x30      ====        or s0, t0, t5
                                                  30'd    11048    : data = 32'h    00BDBB33    ;    //    sltu x22 x27 x11      ====        sltu s6, s11, a1
                                                  30'd    11049    : data = 32'h    414BD393    ;    //    srai x7 x23 20      ====        srai t2, s7, 20
                                                  30'd    11050    : data = 32'h    404D5293    ;    //    srai x5 x26 4      ====        srai t0, s10, 4
                                                  30'd    11051    : data = 32'h    00E00FB3    ;    //    add x31 x0 x14      ====        add t6, zero, a4
                                                  30'd    11052    : data = 32'h    00F85333    ;    //    srl x6 x16 x15      ====        srl t1, a6, a5
                                                  30'd    11053    : data = 32'h    09CF7193    ;    //    andi x3 x30 156      ====        andi gp, t5, 156
                                                  30'd    11054    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11055    : data = 32'h    40425093    ;    //    srai x1 x4 4      ====        srai ra, tp, 4
                                                  30'd    11056    : data = 32'h    40E2D793    ;    //    srai x15 x5 14      ====        srai a5, t0, 14
                                                  30'd    11057    : data = 32'h    41390633    ;    //    sub x12 x18 x19      ====        sub a2, s2, s3
                                                  30'd    11058    : data = 32'h    40BE0A33    ;    //    sub x20 x28 x11      ====        sub s4, t3, a1
                                                  30'd    11059    : data = 32'h    5B2B3093    ;    //    sltiu x1 x22 1458      ====        sltiu ra, s6, 1458
                                                  30'd    11060    : data = 32'h    4014D0B3    ;    //    sra x1 x9 x1      ====        sra ra, s1, ra
                                                  30'd    11061    : data = 32'h    0183B1B3    ;    //    sltu x3 x7 x24      ====        sltu gp, t2, s8
                                                  30'd    11062    : data = 32'h    01BB9993    ;    //    slli x19 x23 27      ====        slli s3, s7, 27
                                                  30'd    11063    : data = 32'h    4198DD13    ;    //    srai x26 x17 25      ====        srai s10, a7, 25
                                                  30'd    11064    : data = 32'h    2D96B397    ;    //    auipc x7 186731      ====        auipc t2, 186731
                                                  30'd    11065    : data = 32'h    0129B2B3    ;    //    sltu x5 x19 x18      ====        sltu t0, s3, s2
                                                  30'd    11066    : data = 32'h    CA112CB7    ;    //    lui x25 827666      ====        lui s9, 827666
                                                  30'd    11067    : data = 32'h    14D8B113    ;    //    sltiu x2 x17 333      ====        sltiu sp, a7, 333
                                                  30'd    11068    : data = 32'h    00A7D493    ;    //    srli x9 x15 10      ====        srli s1, a5, 10
                                                  30'd    11069    : data = 32'h    40130BB3    ;    //    sub x23 x6 x1      ====        sub s7, t1, ra
                                                  30'd    11070    : data = 32'h    009446B3    ;    //    xor x13 x8 x9      ====        xor a3, s0, s1
                                                  30'd    11071    : data = 32'h    7F974B17    ;    //    auipc x22 522612      ====        auipc s6, 522612
                                                  30'd    11072    : data = 32'h    BB5DAF93    ;    //    slti x31 x27 -1099      ====        slti t6, s11, -1099
                                                  30'd    11073    : data = 32'h    00D24B33    ;    //    xor x22 x4 x13      ====        xor s6, tp, a3
                                                  30'd    11074    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11075    : data = 32'h    00A5DE93    ;    //    srli x29 x11 10      ====        srli t4, a1, 10
                                                  30'd    11076    : data = 32'h    5B87BF93    ;    //    sltiu x31 x15 1464      ====        sltiu t6, a5, 1464
                                                  30'd    11077    : data = 32'h    DCE9AB93    ;    //    slti x23 x19 -562      ====        slti s7, s3, -562
                                                  30'd    11078    : data = 32'h    411DD4B3    ;    //    sra x9 x27 x17      ====        sra s1, s11, a7
                                                  30'd    11079    : data = 32'h    CB9978B7    ;    //    lui x17 833943      ====        lui a7, 833943
                                                  30'd    11080    : data = 32'h    0155DA13    ;    //    srli x20 x11 21      ====        srli s4, a1, 21
                                                  30'd    11081    : data = 32'h    4026D413    ;    //    srai x8 x13 2      ====        srai s0, a3, 2
                                                  30'd    11082    : data = 32'h    015A66B3    ;    //    or x13 x20 x21      ====        or a3, s4, s5
                                                  30'd    11083    : data = 32'h    00A11593    ;    //    slli x11 x2 10      ====        slli a1, sp, 10
                                                  30'd    11084    : data = 32'h    DE024613    ;    //    xori x12 x4 -544      ====        xori a2, tp, -544
                                                  30'd    11085    : data = 32'h    B0BA3497    ;    //    auipc x9 723875      ====        auipc s1, 723875
                                                  30'd    11086    : data = 32'h    1A2D4E93    ;    //    xori x29 x26 418      ====        xori t4, s10, 418
                                                  30'd    11087    : data = 32'h    009E98B3    ;    //    sll x17 x29 x9      ====        sll a7, t4, s1
                                                  30'd    11088    : data = 32'h    5CEB2693    ;    //    slti x13 x22 1486      ====        slti a3, s6, 1486
                                                  30'd    11089    : data = 32'h    00959B33    ;    //    sll x22 x11 x9      ====        sll s6, a1, s1
                                                  30'd    11090    : data = 32'h    0137D3B3    ;    //    srl x7 x15 x19      ====        srl t2, a5, s3
                                                  30'd    11091    : data = 32'h    40988933    ;    //    sub x18 x17 x9      ====        sub s2, a7, s1
                                                  30'd    11092    : data = 32'h    8071ED93    ;    //    ori x27 x3 -2041      ====        ori s11, gp, -2041
                                                  30'd    11093    : data = 32'h    41695E33    ;    //    sra x28 x18 x22      ====        sra t3, s2, s6
                                                  30'd    11094    : data = 32'h    069E5897    ;    //    auipc x17 27109      ====        auipc a7, 27109
                                                  30'd    11095    : data = 32'h    AB256B13    ;    //    ori x22 x10 -1358      ====        ori s6, a0, -1358
                                                  30'd    11096    : data = 32'h    006C5733    ;    //    srl x14 x24 x6      ====        srl a4, s8, t1
                                                  30'd    11097    : data = 32'h    403E8733    ;    //    sub x14 x29 x3      ====        sub a4, t4, gp
                                                  30'd    11098    : data = 32'h    00EBB133    ;    //    sltu x2 x23 x14      ====        sltu sp, s7, a4
                                                  30'd    11099    : data = 32'h    00119FB3    ;    //    sll x31 x3 x1      ====        sll t6, gp, ra
                                                  30'd    11100    : data = 32'h    00887E33    ;    //    and x28 x16 x8      ====        and t3, a6, s0
                                                  30'd    11101    : data = 32'h    018DEEB3    ;    //    or x29 x27 x24      ====        or t4, s11, s8
                                                  30'd    11102    : data = 32'h    41B78FB3    ;    //    sub x31 x15 x27      ====        sub t6, a5, s11
                                                  30'd    11103    : data = 32'h    8C00E313    ;    //    ori x6 x1 -1856      ====        ori t1, ra, -1856
                                                  30'd    11104    : data = 32'h    BB564313    ;    //    xori x6 x12 -1099      ====        xori t1, a2, -1099
                                                  30'd    11105    : data = 32'h    01C47033    ;    //    and x0 x8 x28      ====        and zero, s0, t3
                                                  30'd    11106    : data = 32'h    33E64913    ;    //    xori x18 x12 830      ====        xori s2, a2, 830
                                                  30'd    11107    : data = 32'h    BE298093    ;    //    addi x1 x19 -1054      ====        addi ra, s3, -1054
                                                  30'd    11108    : data = 32'h    A51C2113    ;    //    slti x2 x24 -1455      ====        slti sp, s8, -1455
                                                  30'd    11109    : data = 32'h    E23ABC93    ;    //    sltiu x25 x21 -477      ====        sltiu s9, s5, -477
                                                  30'd    11110    : data = 32'h    F893E893    ;    //    ori x17 x7 -119      ====        ori a7, t2, -119
                                                  30'd    11111    : data = 32'h    2906A993    ;    //    slti x19 x13 656      ====        slti s3, a3, 656
                                                  30'd    11112    : data = 32'h    405353B3    ;    //    sra x7 x6 x5      ====        sra t2, t1, t0
                                                  30'd    11113    : data = 32'h    009E1D33    ;    //    sll x26 x28 x9      ====        sll s10, t3, s1
                                                  30'd    11114    : data = 32'h    ADE50F93    ;    //    addi x31 x10 -1314      ====        addi t6, a0, -1314
                                                  30'd    11115    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11116    : data = 32'h    00AA70B3    ;    //    and x1 x20 x10      ====        and ra, s4, a0
                                                  30'd    11117    : data = 32'h    1CECC993    ;    //    xori x19 x25 462      ====        xori s3, s9, 462
                                                  30'd    11118    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11119    : data = 32'h    00C29F93    ;    //    slli x31 x5 12      ====        slli t6, t0, 12
                                                  30'd    11120    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11121    : data = 32'h    0059DDB3    ;    //    srl x27 x19 x5      ====        srl s11, s3, t0
                                                  30'd    11122    : data = 32'h    003D22B3    ;    //    slt x5 x26 x3      ====        slt t0, s10, gp
                                                  30'd    11123    : data = 32'h    2304FA93    ;    //    andi x21 x9 560      ====        andi s5, s1, 560
                                                  30'd    11124    : data = 32'h    01D224B3    ;    //    slt x9 x4 x29      ====        slt s1, tp, t4
                                                  30'd    11125    : data = 32'h    01829C33    ;    //    sll x24 x5 x24      ====        sll s8, t0, s8
                                                  30'd    11126    : data = 32'h    01135E33    ;    //    srl x28 x6 x17      ====        srl t3, t1, a7
                                                  30'd    11127    : data = 32'h    FFCB1497    ;    //    auipc x9 1047729      ====        auipc s1, 1047729
                                                  30'd    11128    : data = 32'h    8DD06937    ;    //    lui x18 580870      ====        lui s2, 580870
                                                  30'd    11129    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11130    : data = 32'h    00021A33    ;    //    sll x20 x4 x0      ====        sll s4, tp, zero
                                                  30'd    11131    : data = 32'h    AC1B4D93    ;    //    xori x27 x22 -1343      ====        xori s11, s6, -1343
                                                  30'd    11132    : data = 32'h    006CE2B3    ;    //    or x5 x25 x6      ====        or t0, s9, t1
                                                  30'd    11133    : data = 32'h    01434DB3    ;    //    xor x27 x6 x20      ====        xor s11, t1, s4
                                                  30'd    11134    : data = 32'h    EA950413    ;    //    addi x8 x10 -343      ====        addi s0, a0, -343
                                                  30'd    11135    : data = 32'h    D0B80293    ;    //    addi x5 x16 -757      ====        addi t0, a6, -757
                                                  30'd    11136    : data = 32'h    09067E93    ;    //    andi x29 x12 144      ====        andi t4, a2, 144
                                                  30'd    11137    : data = 32'h    89BAA937    ;    //    lui x18 564138      ====        lui s2, 564138
                                                  30'd    11138    : data = 32'h    01104633    ;    //    xor x12 x0 x17      ====        xor a2, zero, a7
                                                  30'd    11139    : data = 32'h    0111F833    ;    //    and x16 x3 x17      ====        and a6, gp, a7
                                                  30'd    11140    : data = 32'h    011CCDB3    ;    //    xor x27 x25 x17      ====        xor s11, s9, a7
                                                  30'd    11141    : data = 32'h    4EAB2B13    ;    //    slti x22 x22 1258      ====        slti s6, s6, 1258
                                                  30'd    11142    : data = 32'h    40B18E33    ;    //    sub x28 x3 x11      ====        sub t3, gp, a1
                                                  30'd    11143    : data = 32'h    0183AEB3    ;    //    slt x29 x7 x24      ====        slt t4, t2, s8
                                                  30'd    11144    : data = 32'h    E5AC4693    ;    //    xori x13 x24 -422      ====        xori a3, s8, -422
                                                  30'd    11145    : data = 32'h    40FADD93    ;    //    srai x27 x21 15      ====        srai s11, s5, 15
                                                  30'd    11146    : data = 32'h    00E0BB33    ;    //    sltu x22 x1 x14      ====        sltu s6, ra, a4
                                                  30'd    11147    : data = 32'h    01A3AC33    ;    //    slt x24 x7 x26      ====        slt s8, t2, s10
                                                  30'd    11148    : data = 32'h    40DB5AB3    ;    //    sra x21 x22 x13      ====        sra s5, s6, a3
                                                  30'd    11149    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11150    : data = 32'h    01639093    ;    //    slli x1 x7 22      ====        slli ra, t2, 22
                                                  30'd    11151    : data = 32'h    405CDDB3    ;    //    sra x27 x25 x5      ====        sra s11, s9, t0
                                                  30'd    11152    : data = 32'h    41EB0D33    ;    //    sub x26 x22 x30      ====        sub s10, s6, t5
                                                  30'd    11153    : data = 32'h    007AF5B3    ;    //    and x11 x21 x7      ====        and a1, s5, t2
                                                  30'd    11154    : data = 32'h    E711AD37    ;    //    lui x26 946458      ====        lui s10, 946458
                                                  30'd    11155    : data = 32'h    004FD613    ;    //    srli x12 x31 4      ====        srli a2, t6, 4
                                                  30'd    11156    : data = 32'h    40F90833    ;    //    sub x16 x18 x15      ====        sub a6, s2, a5
                                                  30'd    11157    : data = 32'h    DF600293    ;    //    addi x5 x0 -522      ====        addi t0, zero, -522
                                                  30'd    11158    : data = 32'h    4EF251B7    ;    //    lui x3 323365      ====        lui gp, 323365
                                                  30'd    11159    : data = 32'h    41705E13    ;    //    srai x28 x0 23      ====        srai t3, zero, 23
                                                  30'd    11160    : data = 32'h    7B644193    ;    //    xori x3 x8 1974      ====        xori gp, s0, 1974
                                                  30'd    11161    : data = 32'h    0135A0B3    ;    //    slt x1 x11 x19      ====        slt ra, a1, s3
                                                  30'd    11162    : data = 32'h    B119B313    ;    //    sltiu x6 x19 -1263      ====        sltiu t1, s3, -1263
                                                  30'd    11163    : data = 32'h    407389B3    ;    //    sub x19 x7 x7      ====        sub s3, t2, t2
                                                  30'd    11164    : data = 32'h    00A27333    ;    //    and x6 x4 x10      ====        and t1, tp, a0
                                                  30'd    11165    : data = 32'h    C0D4CD13    ;    //    xori x26 x9 -1011      ====        xori s10, s1, -1011
                                                  30'd    11166    : data = 32'h    8F997393    ;    //    andi x7 x18 -1799      ====        andi t2, s2, -1799
                                                  30'd    11167    : data = 32'h    00744D33    ;    //    xor x26 x8 x7      ====        xor s10, s0, t2
                                                  30'd    11168    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11169    : data = 32'h    0197FB33    ;    //    and x22 x15 x25      ====        and s6, a5, s9
                                                  30'd    11170    : data = 32'h    ABD3AC93    ;    //    slti x25 x7 -1347      ====        slti s9, t2, -1347
                                                  30'd    11171    : data = 32'h    402A85B3    ;    //    sub x11 x21 x2      ====        sub a1, s5, sp
                                                  30'd    11172    : data = 32'h    EF63EA93    ;    //    ori x21 x7 -266      ====        ori s5, t2, -266
                                                  30'd    11173    : data = 32'h    012F6E33    ;    //    or x28 x30 x18      ====        or t3, t5, s2
                                                  30'd    11174    : data = 32'h    F5F28313    ;    //    addi x6 x5 -161      ====        addi t1, t0, -161
                                                  30'd    11175    : data = 32'h    00981113    ;    //    slli x2 x16 9      ====        slli sp, a6, 9
                                                  30'd    11176    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11177    : data = 32'h    409CD9B3    ;    //    sra x19 x25 x9      ====        sra s3, s9, s1
                                                  30'd    11178    : data = 32'h    00000613    ;    //    addi x12 x0 0      ====        li a2, 0x0 #start riscv_int_numeric_corner_stream_12
                                                  30'd    11179    : data = 32'h    00000C13    ;    //    addi x24 x0 0      ====        li s8, 0x0
                                                  30'd    11180    : data = 32'h    FFF00D93    ;    //    addi x27 x0 -1      ====        li s11, 0xffffffff
                                                  30'd    11181    : data = 32'h    00000313    ;    //    addi x6 x0 0      ====        li t1, 0x0
                                                  30'd    11182    : data = 32'h    00000093    ;    //    addi x1 x0 0      ====        li ra, 0x0
                                                  30'd    11183    : data = 32'h    FFF00593    ;    //    addi x11 x0 -1      ====        li a1, 0xffffffff
                                                  30'd    11184    : data = 32'h    80000437    ;    //    lui x8 524288      ====        li s0, 0x80000000
                                                  30'd    11185    : data = 32'h    00040413    ;    //    addi x8 x8 0      ====        li s0, 0x80000000
                                                  30'd    11186    : data = 32'h    FFF00E93    ;    //    addi x29 x0 -1      ====        li t4, 0xffffffff
                                                  30'd    11187    : data = 32'h    0CC59A37    ;    //    lui x20 52313      ====        li s4, 0xcc59027
                                                  30'd    11188    : data = 32'h    027A0A13    ;    //    addi x20 x20 39      ====        li s4, 0xcc59027
                                                  30'd    11189    : data = 32'h    80000AB7    ;    //    lui x21 524288      ====        li s5, 0x80000000
                                                  30'd    11190    : data = 32'h    000A8A93    ;    //    addi x21 x21 0      ====        li s5, 0x80000000
                                                  30'd    11191    : data = 32'h    414E85B3    ;    //    sub x11 x29 x20      ====        sub a1, t4, s4
                                                  30'd    11192    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11193    : data = 32'h    3B0A8093    ;    //    addi x1 x21 944      ====        addi ra, s5, 944
                                                  30'd    11194    : data = 32'h    3F07AC37    ;    //    lui x24 258170      ====        lui s8, 258170
                                                  30'd    11195    : data = 32'h    08EA8613    ;    //    addi x12 x21 142      ====        addi a2, s5, 142
                                                  30'd    11196    : data = 32'h    D31CE0B7    ;    //    lui x1 864718      ====        lui ra, 864718
                                                  30'd    11197    : data = 32'h    FF94B0B7    ;    //    lui x1 1046859      ====        lui ra, 1046859
                                                  30'd    11198    : data = 32'h    4911B617    ;    //    auipc x12 299291      ====        auipc a2, 299291
                                                  30'd    11199    : data = 32'h    29416E97    ;    //    auipc x29 168982      ====        auipc t4, 168982
                                                  30'd    11200    : data = 32'h    40160EB3    ;    //    sub x29 x12 x1      ====        sub t4, a2, ra
                                                  30'd    11201    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11202    : data = 32'h    5B37E0B7    ;    //    lui x1 373630      ====        lui ra, 373630
                                                  30'd    11203    : data = 32'h    FF7E1A97    ;    //    auipc x21 1046497      ====        auipc s5, 1046497
                                                  30'd    11204    : data = 32'h    406600B3    ;    //    sub x1 x12 x6      ====        sub ra, a2, t1
                                                  30'd    11205    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11206    : data = 32'h    40B305B3    ;    //    sub x11 x6 x11      ====        sub a1, t1, a1
                                                  30'd    11207    : data = 32'h    7AEE8093    ;    //    addi x1 x29 1966      ====        addi ra, t4, 1966
                                                  30'd    11208    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11209    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11210    : data = 32'h    0BAE8613    ;    //    addi x12 x29 186      ====        addi a2, t4, 186
                                                  30'd    11211    : data = 32'h    01D08C33    ;    //    add x24 x1 x29      ====        add s8, ra, t4
                                                  30'd    11212    : data = 32'h    96FED337    ;    //    lui x6 618477      ====        lui t1, 618477
                                                  30'd    11213    : data = 32'h    01B305B3    ;    //    add x11 x6 x27      ====        add a1, t1, s11
                                                  30'd    11214    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11215    : data = 32'h    00658EB3    ;    //    add x29 x11 x6      ====        add t4, a1, t1
                                                  30'd    11216    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11217    : data = 32'h    024E1337    ;    //    lui x6 9441      ====        lui t1, 9441
                                                  30'd    11218    : data = 32'h    008D85B3    ;    //    add x11 x27 x8      ====        add a1, s11, s0
                                                  30'd    11219    : data = 32'h    00CD80B3    ;    //    add x1 x27 x12      ====        add ra, s11, a2
                                                  30'd    11220    : data = 32'h    798000EF    ;    //    jal x1 1944      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_12
                                                  30'd    11221    : data = 32'h    00B2D593    ;    //    srli x11 x5 11      ====        srli a1, t0, 11
                                                  30'd    11222    : data = 32'h    008F0733    ;    //    add x14 x30 x8      ====        add a4, t5, s0
                                                  30'd    11223    : data = 32'h    092CBE13    ;    //    sltiu x28 x25 146      ====        sltiu t3, s9, 146
                                                  30'd    11224    : data = 32'h    400AD793    ;    //    srai x15 x21 0      ====        srai a5, s5, 0
                                                  30'd    11225    : data = 32'h    416889B3    ;    //    sub x19 x17 x22      ====        sub s3, a7, s6
                                                  30'd    11226    : data = 32'h    017CE2B3    ;    //    or x5 x25 x23      ====        or t0, s9, s7
                                                  30'd    11227    : data = 32'h    01984833    ;    //    xor x16 x16 x25      ====        xor a6, a6, s9
                                                  30'd    11228    : data = 32'h    41C55D33    ;    //    sra x26 x10 x28      ====        sra s10, a0, t3
                                                  30'd    11229    : data = 32'h    01195C93    ;    //    srli x25 x18 17      ====        srli s9, s2, 17
                                                  30'd    11230    : data = 32'h    007F20B3    ;    //    slt x1 x30 x7      ====        slt ra, t5, t2
                                                  30'd    11231    : data = 32'h    27AAF093    ;    //    andi x1 x21 634      ====        andi ra, s5, 634
                                                  30'd    11232    : data = 32'h    01B774B3    ;    //    and x9 x14 x27      ====        and s1, a4, s11
                                                  30'd    11233    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11234    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11235    : data = 32'h    40E10633    ;    //    sub x12 x2 x14      ====        sub a2, sp, a4
                                                  30'd    11236    : data = 32'h    019D9B13    ;    //    slli x22 x27 25      ====        slli s6, s11, 25
                                                  30'd    11237    : data = 32'h    103CFB93    ;    //    andi x23 x25 259      ====        andi s7, s9, 259
                                                  30'd    11238    : data = 32'h    C4258313    ;    //    addi x6 x11 -958      ====        addi t1, a1, -958
                                                  30'd    11239    : data = 32'h    001D8333    ;    //    add x6 x27 x1      ====        add t1, s11, ra
                                                  30'd    11240    : data = 32'h    407205B3    ;    //    sub x11 x4 x7      ====        sub a1, tp, t2
                                                  30'd    11241    : data = 32'h    01F80DB3    ;    //    add x27 x16 x31      ====        add s11, a6, t6
                                                  30'd    11242    : data = 32'h    00C33E33    ;    //    sltu x28 x6 x12      ====        sltu t3, t1, a2
                                                  30'd    11243    : data = 32'h    40518333    ;    //    sub x6 x3 x5      ====        sub t1, gp, t0
                                                  30'd    11244    : data = 32'h    01316DB3    ;    //    or x27 x2 x19      ====        or s11, sp, s3
                                                  30'd    11245    : data = 32'h    00DA34B3    ;    //    sltu x9 x20 x13      ====        sltu s1, s4, a3
                                                  30'd    11246    : data = 32'h    D5FC45B7    ;    //    lui x11 876484      ====        lui a1, 876484
                                                  30'd    11247    : data = 32'h    01D761B3    ;    //    or x3 x14 x29      ====        or gp, a4, t4
                                                  30'd    11248    : data = 32'h    0148A333    ;    //    slt x6 x17 x20      ====        slt t1, a7, s4
                                                  30'd    11249    : data = 32'h    01CFD193    ;    //    srli x3 x31 28      ====        srli gp, t6, 28
                                                  30'd    11250    : data = 32'h    AD011297    ;    //    auipc x5 708625      ====        auipc t0, 708625
                                                  30'd    11251    : data = 32'h    719A2613    ;    //    slti x12 x20 1817      ====        slti a2, s4, 1817
                                                  30'd    11252    : data = 32'h    009209B3    ;    //    add x19 x4 x9      ====        add s3, tp, s1
                                                  30'd    11253    : data = 32'h    D59BF693    ;    //    andi x13 x23 -679      ====        andi a3, s7, -679
                                                  30'd    11254    : data = 32'h    632D6A97    ;    //    auipc x21 406230      ====        auipc s5, 406230
                                                  30'd    11255    : data = 32'h    01A65433    ;    //    srl x8 x12 x26      ====        srl s0, a2, s10
                                                  30'd    11256    : data = 32'h    00F2BE33    ;    //    sltu x28 x5 x15      ====        sltu t3, t0, a5
                                                  30'd    11257    : data = 32'h    00239993    ;    //    slli x19 x7 2      ====        slli s3, t2, 2
                                                  30'd    11258    : data = 32'h    01D624B3    ;    //    slt x9 x12 x29      ====        slt s1, a2, t4
                                                  30'd    11259    : data = 32'h    00C75733    ;    //    srl x14 x14 x12      ====        srl a4, a4, a2
                                                  30'd    11260    : data = 32'h    38C93B93    ;    //    sltiu x23 x18 908      ====        sltiu s7, s2, 908
                                                  30'd    11261    : data = 32'h    3F0F2713    ;    //    slti x14 x30 1008      ====        slti a4, t5, 1008
                                                  30'd    11262    : data = 32'h    41E15BB3    ;    //    sra x23 x2 x30      ====        sra s7, sp, t5
                                                  30'd    11263    : data = 32'h    016C2BB3    ;    //    slt x23 x24 x22      ====        slt s7, s8, s6
                                                  30'd    11264    : data = 32'h    A1C9EE93    ;    //    ori x29 x19 -1508      ====        ori t4, s3, -1508
                                                  30'd    11265    : data = 32'h    0197BFB3    ;    //    sltu x31 x15 x25      ====        sltu t6, a5, s9
                                                  30'd    11266    : data = 32'h    41045B93    ;    //    srai x23 x8 16      ====        srai s7, s0, 16
                                                  30'd    11267    : data = 32'h    AF0D6D13    ;    //    ori x26 x26 -1296      ====        ori s10, s10, -1296
                                                  30'd    11268    : data = 32'h    39ACFB13    ;    //    andi x22 x25 922      ====        andi s6, s9, 922
                                                  30'd    11269    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11270    : data = 32'h    01A927B3    ;    //    slt x15 x18 x26      ====        slt a5, s2, s10
                                                  30'd    11271    : data = 32'h    0194FFB3    ;    //    and x31 x9 x25      ====        and t6, s1, s9
                                                  30'd    11272    : data = 32'h    00D85BB3    ;    //    srl x23 x16 x13      ====        srl s7, a6, a3
                                                  30'd    11273    : data = 32'h    E58CFC17    ;    //    auipc x24 940239      ====        auipc s8, 940239
                                                  30'd    11274    : data = 32'h    00085013    ;    //    srli x0 x16 0      ====        srli zero, a6, 0
                                                  30'd    11275    : data = 32'h    AEF5CC93    ;    //    xori x25 x11 -1297      ====        xori s9, a1, -1297
                                                  30'd    11276    : data = 32'h    8AF42313    ;    //    slti x6 x8 -1873      ====        slti t1, s0, -1873
                                                  30'd    11277    : data = 32'h    00283C33    ;    //    sltu x24 x16 x2      ====        sltu s8, a6, sp
                                                  30'd    11278    : data = 32'h    0015E5B3    ;    //    or x11 x11 x1      ====        or a1, a1, ra
                                                  30'd    11279    : data = 32'h    01740D33    ;    //    add x26 x8 x23      ====        add s10, s0, s7
                                                  30'd    11280    : data = 32'h    018432B3    ;    //    sltu x5 x8 x24      ====        sltu t0, s0, s8
                                                  30'd    11281    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11282    : data = 32'h    415D53B3    ;    //    sra x7 x26 x21      ====        sra t2, s10, s5
                                                  30'd    11283    : data = 32'h    01FD4FB3    ;    //    xor x31 x26 x31      ====        xor t6, s10, t6
                                                  30'd    11284    : data = 32'h    01A81833    ;    //    sll x16 x16 x26      ====        sll a6, a6, s10
                                                  30'd    11285    : data = 32'h    011D5CB3    ;    //    srl x25 x26 x17      ====        srl s9, s10, a7
                                                  30'd    11286    : data = 32'h    403B5CB3    ;    //    sra x25 x22 x3      ====        sra s9, s6, gp
                                                  30'd    11287    : data = 32'h    8BEFD717    ;    //    auipc x14 573181      ====        auipc a4, 573181
                                                  30'd    11288    : data = 32'h    0015CCB3    ;    //    xor x25 x11 x1      ====        xor s9, a1, ra
                                                  30'd    11289    : data = 32'h    F0F2C293    ;    //    xori x5 x5 -241      ====        xori t0, t0, -241
                                                  30'd    11290    : data = 32'h    6E7D7113    ;    //    andi x2 x26 1767      ====        andi sp, s10, 1767
                                                  30'd    11291    : data = 32'h    01226633    ;    //    or x12 x4 x18      ====        or a2, tp, s2
                                                  30'd    11292    : data = 32'h    001E1713    ;    //    slli x14 x28 1      ====        slli a4, t3, 1
                                                  30'd    11293    : data = 32'h    504F8713    ;    //    addi x14 x31 1284      ====        addi a4, t6, 1284
                                                  30'd    11294    : data = 32'h    075A7793    ;    //    andi x15 x20 117      ====        andi a5, s4, 117
                                                  30'd    11295    : data = 32'h    006BBB33    ;    //    sltu x22 x23 x6      ====        sltu s6, s7, t1
                                                  30'd    11296    : data = 32'h    AC168313    ;    //    addi x6 x13 -1343      ====        addi t1, a3, -1343
                                                  30'd    11297    : data = 32'h    4173D713    ;    //    srai x14 x7 23      ====        srai a4, t2, 23
                                                  30'd    11298    : data = 32'h    3F6C5097    ;    //    auipc x1 259781      ====        auipc ra, 259781
                                                  30'd    11299    : data = 32'h    01741733    ;    //    sll x14 x8 x23      ====        sll a4, s0, s7
                                                  30'd    11300    : data = 32'h    B4BC0317    ;    //    auipc x6 740288      ====        auipc t1, 740288
                                                  30'd    11301    : data = 32'h    E3F72793    ;    //    slti x15 x14 -449      ====        slti a5, a4, -449
                                                  30'd    11302    : data = 32'h    00741713    ;    //    slli x14 x8 7      ====        slli a4, s0, 7
                                                  30'd    11303    : data = 32'h    512E4493    ;    //    xori x9 x28 1298      ====        xori s1, t3, 1298
                                                  30'd    11304    : data = 32'h    41828B33    ;    //    sub x22 x5 x24      ====        sub s6, t0, s8
                                                  30'd    11305    : data = 32'h    00EFA4B3    ;    //    slt x9 x31 x14      ====        slt s1, t6, a4
                                                  30'd    11306    : data = 32'h    0037D133    ;    //    srl x2 x15 x3      ====        srl sp, a5, gp
                                                  30'd    11307    : data = 32'h    19F7AA13    ;    //    slti x20 x15 415      ====        slti s4, a5, 415
                                                  30'd    11308    : data = 32'h    05F17E13    ;    //    andi x28 x2 95      ====        andi t3, sp, 95
                                                  30'd    11309    : data = 32'h    01CBE333    ;    //    or x6 x23 x28      ====        or t1, s7, t3
                                                  30'd    11310    : data = 32'h    41465D13    ;    //    srai x26 x12 20      ====        srai s10, a2, 20
                                                  30'd    11311    : data = 32'h    40195E13    ;    //    srai x28 x18 1      ====        srai t3, s2, 1
                                                  30'd    11312    : data = 32'h    2C033A13    ;    //    sltiu x20 x6 704      ====        sltiu s4, t1, 704
                                                  30'd    11313    : data = 32'h    00209413    ;    //    slli x8 x1 2      ====        slli s0, ra, 2
                                                  30'd    11314    : data = 32'h    005C28B3    ;    //    slt x17 x24 x5      ====        slt a7, s8, t0
                                                  30'd    11315    : data = 32'h    37277593    ;    //    andi x11 x14 882      ====        andi a1, a4, 882
                                                  30'd    11316    : data = 32'h    A0750B37    ;    //    lui x22 657232      ====        lui s6, 657232
                                                  30'd    11317    : data = 32'h    007AC933    ;    //    xor x18 x21 x7      ====        xor s2, s5, t2
                                                  30'd    11318    : data = 32'h    0195ED33    ;    //    or x26 x11 x25      ====        or s10, a1, s9
                                                  30'd    11319    : data = 32'h    407C5F93    ;    //    srai x31 x24 7      ====        srai t6, s8, 7
                                                  30'd    11320    : data = 32'h    95E34793    ;    //    xori x15 x6 -1698      ====        xori a5, t1, -1698
                                                  30'd    11321    : data = 32'h    0DCE7E13    ;    //    andi x28 x28 220      ====        andi t3, t3, 220
                                                  30'd    11322    : data = 32'h    41365E93    ;    //    srai x29 x12 19      ====        srai t4, a2, 19
                                                  30'd    11323    : data = 32'h    01F85613    ;    //    srli x12 x16 31      ====        srli a2, a6, 31
                                                  30'd    11324    : data = 32'h    00391033    ;    //    sll x0 x18 x3      ====        sll zero, s2, gp
                                                  30'd    11325    : data = 32'h    403C5B33    ;    //    sra x22 x24 x3      ====        sra s6, s8, gp
                                                  30'd    11326    : data = 32'h    B1020E13    ;    //    addi x28 x4 -1264      ====        addi t3, tp, -1264
                                                  30'd    11327    : data = 32'h    40CA80B3    ;    //    sub x1 x21 x12      ====        sub ra, s5, a2
                                                  30'd    11328    : data = 32'h    013E2733    ;    //    slt x14 x28 x19      ====        slt a4, t3, s3
                                                  30'd    11329    : data = 32'h    00C58033    ;    //    add x0 x11 x12      ====        add zero, a1, a2
                                                  30'd    11330    : data = 32'h    B3657913    ;    //    andi x18 x10 -1226      ====        andi s2, a0, -1226
                                                  30'd    11331    : data = 32'h    00000B13    ;    //    addi x22 x0 0      ====        li s6, 0x0 #start riscv_int_numeric_corner_stream_0
                                                  30'd    11332    : data = 32'h    953AB9B7    ;    //    lui x19 611243      ====        li s3, 0x953aaa71
                                                  30'd    11333    : data = 32'h    A7198993    ;    //    addi x19 x19 -1423      ====        li s3, 0x953aaa71
                                                  30'd    11334    : data = 32'h    FFF00E93    ;    //    addi x29 x0 -1      ====        li t4, 0xffffffff
                                                  30'd    11335    : data = 32'h    00000B93    ;    //    addi x23 x0 0      ====        li s7, 0x0
                                                  30'd    11336    : data = 32'h    800008B7    ;    //    lui x17 524288      ====        li a7, 0x80000000
                                                  30'd    11337    : data = 32'h    00088893    ;    //    addi x17 x17 0      ====        li a7, 0x80000000
                                                  30'd    11338    : data = 32'h    FFF00713    ;    //    addi x14 x0 -1      ====        li a4, 0xffffffff
                                                  30'd    11339    : data = 32'h    FFF00193    ;    //    addi x3 x0 -1      ====        li gp, 0xffffffff
                                                  30'd    11340    : data = 32'h    FFF00413    ;    //    addi x8 x0 -1      ====        li s0, 0xffffffff
                                                  30'd    11341    : data = 32'h    FFF00D93    ;    //    addi x27 x0 -1      ====        li s11, 0xffffffff
                                                  30'd    11342    : data = 32'h    80000D37    ;    //    lui x26 524288      ====        li s10, 0x80000000
                                                  30'd    11343    : data = 32'h    000D0D13    ;    //    addi x26 x26 0      ====        li s10, 0x80000000
                                                  30'd    11344    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11345    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11346    : data = 32'h    00888733    ;    //    add x14 x17 x8      ====        add a4, a7, s0
                                                  30'd    11347    : data = 32'h    413D8733    ;    //    sub x14 x27 x19      ====        sub a4, s11, s3
                                                  30'd    11348    : data = 32'h    76925E97    ;    //    auipc x29 485669      ====        auipc t4, 485669
                                                  30'd    11349    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11350    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11351    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11352    : data = 32'h    00EB09B3    ;    //    add x19 x22 x14      ====        add s3, s6, a4
                                                  30'd    11353    : data = 32'h    4EE03B17    ;    //    auipc x22 323075      ====        auipc s6, 323075
                                                  30'd    11354    : data = 32'h    923B3EB7    ;    //    lui x29 598963      ====        lui t4, 598963
                                                  30'd    11355    : data = 32'h    15D42B17    ;    //    auipc x22 89410      ====        auipc s6, 89410
                                                  30'd    11356    : data = 32'h    003D88B3    ;    //    add x17 x27 x3      ====        add a7, s11, gp
                                                  30'd    11357    : data = 32'h    EDACAB37    ;    //    lui x22 973514      ====        lui s6, 973514
                                                  30'd    11358    : data = 32'h    C036F737    ;    //    lui x14 787311      ====        lui a4, 787311
                                                  30'd    11359    : data = 32'h    016E8BB3    ;    //    add x23 x29 x22      ====        add s7, t4, s6
                                                  30'd    11360    : data = 32'h    5EED0B93    ;    //    addi x23 x26 1518      ====        addi s7, s10, 1518
                                                  30'd    11361    : data = 32'h    D76EB897    ;    //    auipc x17 882411      ====        auipc a7, 882411
                                                  30'd    11362    : data = 32'h    01640B33    ;    //    add x22 x8 x22      ====        add s6, s0, s6
                                                  30'd    11363    : data = 32'h    E7309B37    ;    //    lui x22 946953      ====        lui s6, 946953
                                                  30'd    11364    : data = 32'h    E4598193    ;    //    addi x3 x19 -443      ====        addi gp, s3, -443
                                                  30'd    11365    : data = 32'h    1DDB0893    ;    //    addi x17 x22 477      ====        addi a7, s6, 477
                                                  30'd    11366    : data = 32'h    936721B7    ;    //    lui x3 603762      ====        lui gp, 603762
                                                  30'd    11367    : data = 32'h    54C000EF    ;    //    jal x1 1356      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_0
                                                  30'd    11368    : data = 32'h    7BED4913    ;    //    xori x18 x26 1982      ====        xori s2, s10, 1982
                                                  30'd    11369    : data = 32'h    004E5D93    ;    //    srli x27 x28 4      ====        srli s11, t3, 4
                                                  30'd    11370    : data = 32'h    01A3C6B3    ;    //    xor x13 x7 x26      ====        xor a3, t2, s10
                                                  30'd    11371    : data = 32'h    B3C17C13    ;    //    andi x24 x2 -1220      ====        andi s8, sp, -1220
                                                  30'd    11372    : data = 32'h    003C9193    ;    //    slli x3 x25 3      ====        slli gp, s9, 3
                                                  30'd    11373    : data = 32'h    0174CAB3    ;    //    xor x21 x9 x23      ====        xor s5, s1, s7
                                                  30'd    11374    : data = 32'h    004D06B3    ;    //    add x13 x26 x4      ====        add a3, s10, tp
                                                  30'd    11375    : data = 32'h    419EDD93    ;    //    srai x27 x29 25      ====        srai s11, t4, 25
                                                  30'd    11376    : data = 32'h    409ED713    ;    //    srai x14 x29 9      ====        srai a4, t4, 9
                                                  30'd    11377    : data = 32'h    010C2D33    ;    //    slt x26 x24 x16      ====        slt s10, s8, a6
                                                  30'd    11378    : data = 32'h    01ECD2B3    ;    //    srl x5 x25 x30      ====        srl t0, s9, t5
                                                  30'd    11379    : data = 32'h    007953B3    ;    //    srl x7 x18 x7      ====        srl t2, s2, t2
                                                  30'd    11380    : data = 32'h    419CD433    ;    //    sra x8 x25 x25      ====        sra s0, s9, s9
                                                  30'd    11381    : data = 32'h    00FCF4B3    ;    //    and x9 x25 x15      ====        and s1, s9, a5
                                                  30'd    11382    : data = 32'h    007A3CB3    ;    //    sltu x25 x20 x7      ====        sltu s9, s4, t2
                                                  30'd    11383    : data = 32'h    004F8BB3    ;    //    add x23 x31 x4      ====        add s7, t6, tp
                                                  30'd    11384    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11385    : data = 32'h    01450033    ;    //    add x0 x10 x20      ====        add zero, a0, s4
                                                  30'd    11386    : data = 32'h    8337C693    ;    //    xori x13 x15 -1997      ====        xori a3, a5, -1997
                                                  30'd    11387    : data = 32'h    004D7DB3    ;    //    and x27 x26 x4      ====        and s11, s10, tp
                                                  30'd    11388    : data = 32'h    5D6EBA93    ;    //    sltiu x21 x29 1494      ====        sltiu s5, t4, 1494
                                                  30'd    11389    : data = 32'h    BF46F393    ;    //    andi x7 x13 -1036      ====        andi t2, a3, -1036
                                                  30'd    11390    : data = 32'h    9160E013    ;    //    ori x0 x1 -1770      ====        ori zero, ra, -1770
                                                  30'd    11391    : data = 32'h    01273BB3    ;    //    sltu x23 x14 x18      ====        sltu s7, a4, s2
                                                  30'd    11392    : data = 32'h    701D6E13    ;    //    ori x28 x26 1793      ====        ori t3, s10, 1793
                                                  30'd    11393    : data = 32'h    0023C633    ;    //    xor x12 x7 x2      ====        xor a2, t2, sp
                                                  30'd    11394    : data = 32'h    41EEDC93    ;    //    srai x25 x29 30      ====        srai s9, t4, 30
                                                  30'd    11395    : data = 32'h    41EE8FB3    ;    //    sub x31 x29 x30      ====        sub t6, t4, t5
                                                  30'd    11396    : data = 32'h    457DCE37    ;    //    lui x28 284636      ====        lui t3, 284636
                                                  30'd    11397    : data = 32'h    CC8EE437    ;    //    lui x8 837870      ====        lui s0, 837870
                                                  30'd    11398    : data = 32'h    008D7CB3    ;    //    and x25 x26 x8      ====        and s9, s10, s0
                                                  30'd    11399    : data = 32'h    04928713    ;    //    addi x14 x5 73      ====        addi a4, t0, 73
                                                  30'd    11400    : data = 32'h    5EE4C813    ;    //    xori x16 x9 1518      ====        xori a6, s1, 1518
                                                  30'd    11401    : data = 32'h    E8BB8393    ;    //    addi x7 x23 -373      ====        addi t2, s7, -373
                                                  30'd    11402    : data = 32'h    00E783B3    ;    //    add x7 x15 x14      ====        add t2, a5, a4
                                                  30'd    11403    : data = 32'h    00E85A13    ;    //    srli x20 x16 14      ====        srli s4, a6, 14
                                                  30'd    11404    : data = 32'h    00469333    ;    //    sll x6 x13 x4      ====        sll t1, a3, tp
                                                  30'd    11405    : data = 32'h    418DD613    ;    //    srai x12 x27 24      ====        srai a2, s11, 24
                                                  30'd    11406    : data = 32'h    005DEEB3    ;    //    or x29 x27 x5      ====        or t4, s11, t0
                                                  30'd    11407    : data = 32'h    0DCCB593    ;    //    sltiu x11 x25 220      ====        sltiu a1, s9, 220
                                                  30'd    11408    : data = 32'h    003990B3    ;    //    sll x1 x19 x3      ====        sll ra, s3, gp
                                                  30'd    11409    : data = 32'h    BB4F0093    ;    //    addi x1 x30 -1100      ====        addi ra, t5, -1100
                                                  30'd    11410    : data = 32'h    002750B3    ;    //    srl x1 x14 x2      ====        srl ra, a4, sp
                                                  30'd    11411    : data = 32'h    87B1F193    ;    //    andi x3 x3 -1925      ====        andi gp, gp, -1925
                                                  30'd    11412    : data = 32'h    67F3C493    ;    //    xori x9 x7 1663      ====        xori s1, t2, 1663
                                                  30'd    11413    : data = 32'h    40C8D7B3    ;    //    sra x15 x17 x12      ====        sra a5, a7, a2
                                                  30'd    11414    : data = 32'h    41065313    ;    //    srai x6 x12 16      ====        srai t1, a2, 16
                                                  30'd    11415    : data = 32'h    F9C63893    ;    //    sltiu x17 x12 -100      ====        sltiu a7, a2, -100
                                                  30'd    11416    : data = 32'h    FD524313    ;    //    xori x6 x4 -43      ====        xori t1, tp, -43
                                                  30'd    11417    : data = 32'h    AB7EE893    ;    //    ori x17 x29 -1353      ====        ori a7, t4, -1353
                                                  30'd    11418    : data = 32'h    00D862B3    ;    //    or x5 x16 x13      ====        or t0, a6, a3
                                                  30'd    11419    : data = 32'h    AD098093    ;    //    addi x1 x19 -1328      ====        addi ra, s3, -1328
                                                  30'd    11420    : data = 32'h    A8E66193    ;    //    ori x3 x12 -1394      ====        ori gp, a2, -1394
                                                  30'd    11421    : data = 32'h    AF93BB93    ;    //    sltiu x23 x7 -1287      ====        sltiu s7, t2, -1287
                                                  30'd    11422    : data = 32'h    8517C093    ;    //    xori x1 x15 -1967      ====        xori ra, a5, -1967
                                                  30'd    11423    : data = 32'h    B30C19B7    ;    //    lui x19 733377      ====        lui s3, 733377
                                                  30'd    11424    : data = 32'h    01837FB3    ;    //    and x31 x6 x24      ====        and t6, t1, s8
                                                  30'd    11425    : data = 32'h    002D5B33    ;    //    srl x22 x26 x2      ====        srl s6, s10, sp
                                                  30'd    11426    : data = 32'h    E470CB93    ;    //    xori x23 x1 -441      ====        xori s7, ra, -441
                                                  30'd    11427    : data = 32'h    B7E0C113    ;    //    xori x2 x1 -1154      ====        xori sp, ra, -1154
                                                  30'd    11428    : data = 32'h    01DC0733    ;    //    add x14 x24 x29      ====        add a4, s8, t4
                                                  30'd    11429    : data = 32'h    00E1BB33    ;    //    sltu x22 x3 x14      ====        sltu s6, gp, a4
                                                  30'd    11430    : data = 32'h    4181DB33    ;    //    sra x22 x3 x24      ====        sra s6, gp, s8
                                                  30'd    11431    : data = 32'h    00FEC0B3    ;    //    xor x1 x29 x15      ====        xor ra, t4, a5
                                                  30'd    11432    : data = 32'h    016A88B3    ;    //    add x17 x21 x22      ====        add a7, s5, s6
                                                  30'd    11433    : data = 32'h    CAC95B37    ;    //    lui x22 830613      ====        lui s6, 830613
                                                  30'd    11434    : data = 32'h    006BB633    ;    //    sltu x12 x23 x6      ====        sltu a2, s7, t1
                                                  30'd    11435    : data = 32'h    6A557B93    ;    //    andi x23 x10 1701      ====        andi s7, a0, 1701
                                                  30'd    11436    : data = 32'h    40070A33    ;    //    sub x20 x14 x0      ====        sub s4, a4, zero
                                                  30'd    11437    : data = 32'h    00D5F5B3    ;    //    and x11 x11 x13      ====        and a1, a1, a3
                                                  30'd    11438    : data = 32'h    ED13EA13    ;    //    ori x20 x7 -303      ====        ori s4, t2, -303
                                                  30'd    11439    : data = 32'h    416F5B93    ;    //    srai x23 x30 22      ====        srai s7, t5, 22
                                                  30'd    11440    : data = 32'h    00A28933    ;    //    add x18 x5 x10      ====        add s2, t0, a0
                                                  30'd    11441    : data = 32'h    01D86D33    ;    //    or x26 x16 x29      ====        or s10, a6, t4
                                                  30'd    11442    : data = 32'h    29007413    ;    //    andi x8 x0 656      ====        andi s0, zero, 656
                                                  30'd    11443    : data = 32'h    C4A27C13    ;    //    andi x24 x4 -950      ====        andi s8, tp, -950
                                                  30'd    11444    : data = 32'h    01A377B3    ;    //    and x15 x6 x26      ====        and a5, t1, s10
                                                  30'd    11445    : data = 32'h    01D85093    ;    //    srli x1 x16 29      ====        srli ra, a6, 29
                                                  30'd    11446    : data = 32'h    40B60893    ;    //    addi x17 x12 1035      ====        addi a7, a2, 1035
                                                  30'd    11447    : data = 32'h    016A1433    ;    //    sll x8 x20 x22      ====        sll s0, s4, s6
                                                  30'd    11448    : data = 32'h    DDA70113    ;    //    addi x2 x14 -550      ====        addi sp, a4, -550
                                                  30'd    11449    : data = 32'h    00B301B3    ;    //    add x3 x6 x11      ====        add gp, t1, a1
                                                  30'd    11450    : data = 32'h    FAEAFD13    ;    //    andi x26 x21 -82      ====        andi s10, s5, -82
                                                  30'd    11451    : data = 32'h    011E6333    ;    //    or x6 x28 x17      ====        or t1, t3, a7
                                                  30'd    11452    : data = 32'h    C4F53713    ;    //    sltiu x14 x10 -945      ====        sltiu a4, a0, -945
                                                  30'd    11453    : data = 32'h    00AB2BB3    ;    //    slt x23 x22 x10      ====        slt s7, s6, a0
                                                  30'd    11454    : data = 32'h    59D057B7    ;    //    lui x15 367877      ====        lui a5, 367877
                                                  30'd    11455    : data = 32'h    3917E113    ;    //    ori x2 x15 913      ====        ori sp, a5, 913
                                                  30'd    11456    : data = 32'h    003426B3    ;    //    slt x13 x8 x3      ====        slt a3, s0, gp
                                                  30'd    11457    : data = 32'h    0138D633    ;    //    srl x12 x17 x19      ====        srl a2, a7, s3
                                                  30'd    11458    : data = 32'h    40235C33    ;    //    sra x24 x6 x2      ====        sra s8, t1, sp
                                                  30'd    11459    : data = 32'h    0083AE33    ;    //    slt x28 x7 x8      ====        slt t3, t2, s0
                                                  30'd    11460    : data = 32'h    21B0A313    ;    //    slti x6 x1 539      ====        slti t1, ra, 539
                                                  30'd    11461    : data = 32'h    58497593    ;    //    andi x11 x18 1412      ====        andi a1, s2, 1412
                                                  30'd    11462    : data = 32'h    01459633    ;    //    sll x12 x11 x20      ====        sll a2, a1, s4
                                                  30'd    11463    : data = 32'h    12AA2493    ;    //    slti x9 x20 298      ====        slti s1, s4, 298
                                                  30'd    11464    : data = 32'h    AD624713    ;    //    xori x14 x4 -1322      ====        xori a4, tp, -1322
                                                  30'd    11465    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11466    : data = 32'h    0064FD33    ;    //    and x26 x9 x6      ====        and s10, s1, t1
                                                  30'd    11467    : data = 32'h    9C743193    ;    //    sltiu x3 x8 -1593      ====        sltiu gp, s0, -1593
                                                  30'd    11468    : data = 32'h    01379933    ;    //    sll x18 x15 x19      ====        sll s2, a5, s3
                                                  30'd    11469    : data = 32'h    B36CC713    ;    //    xori x14 x25 -1226      ====        xori a4, s9, -1226
                                                  30'd    11470    : data = 32'h    00150E33    ;    //    add x28 x10 x1      ====        add t3, a0, ra
                                                  30'd    11471    : data = 32'h    8A047D13    ;    //    andi x26 x8 -1888      ====        andi s10, s0, -1888
                                                  30'd    11472    : data = 32'h    40E90933    ;    //    sub x18 x18 x14      ====        sub s2, s2, a4
                                                  30'd    11473    : data = 32'h    00553933    ;    //    sltu x18 x10 x5      ====        sltu s2, a0, t0
                                                  30'd    11474    : data = 32'h    B34139B7    ;    //    lui x19 734227      ====        lui s3, 734227
                                                  30'd    11475    : data = 32'h    4084D113    ;    //    srai x2 x9 8      ====        srai sp, s1, 8
                                                  30'd    11476    : data = 32'h    00A4F9B3    ;    //    and x19 x9 x10      ====        and s3, s1, a0
                                                  30'd    11477    : data = 32'h    729A0B37    ;    //    lui x22 469408      ====        lui s6, 469408
                                                  30'd    11478    : data = 32'h    2416BD93    ;    //    sltiu x27 x13 577      ====        sltiu s11, a3, 577
                                                  30'd    11479    : data = 32'h    41A4DA13    ;    //    srai x20 x9 26      ====        srai s4, s1, 26
                                                  30'd    11480    : data = 32'h    01402AB3    ;    //    slt x21 x0 x20      ====        slt s5, zero, s4
                                                  30'd    11481    : data = 32'h    00D25193    ;    //    srli x3 x4 13      ====        srli gp, tp, 13
                                                  30'd    11482    : data = 32'h    00C457B3    ;    //    srl x15 x8 x12      ====        srl a5, s0, a2
                                                  30'd    11483    : data = 32'h    6A490CB7    ;    //    lui x25 435344      ====        lui s9, 435344
                                                  30'd    11484    : data = 32'h    003CACB3    ;    //    slt x25 x25 x3      ====        slt s9, s9, gp
                                                  30'd    11485    : data = 32'h    E6E0DBB7    ;    //    lui x23 945677      ====        lui s7, 945677
                                                  30'd    11486    : data = 32'h    197AD617    ;    //    auipc x12 104365      ====        auipc a2, 104365
                                                  30'd    11487    : data = 32'h    000EE333    ;    //    or x6 x29 x0      ====        or t1, t4, zero
                                                  30'd    11488    : data = 32'h    019A1E13    ;    //    slli x28 x20 25      ====        slli t3, s4, 25
                                                  30'd    11489    : data = 32'h    0A443437    ;    //    lui x8 42051      ====        lui s0, 42051
                                                  30'd    11490    : data = 32'h    014AC8B3    ;    //    xor x17 x21 x20      ====        xor a7, s5, s4
                                                  30'd    11491    : data = 32'h    DA4F6013    ;    //    ori x0 x30 -604      ====        ori zero, t5, -604
                                                  30'd    11492    : data = 32'h    01DCCB33    ;    //    xor x22 x25 x29      ====        xor s6, s9, t4
                                                  30'd    11493    : data = 32'h    8D6EB9B7    ;    //    lui x19 579307      ====        lui s3, 579307
                                                  30'd    11494    : data = 32'h    01D81D13    ;    //    slli x26 x16 29      ====        slli s10, a6, 29
                                                  30'd    11495    : data = 32'h    4BB63393    ;    //    sltiu x7 x12 1211      ====        sltiu t2, a2, 1211
                                                  30'd    11496    : data = 32'h    01C1AD33    ;    //    slt x26 x3 x28      ====        slt s10, gp, t3
                                                  30'd    11497    : data = 32'h    40AFDAB3    ;    //    sra x21 x31 x10      ====        sra s5, t6, a0
                                                  30'd    11498    : data = 32'h    00AAEFB3    ;    //    or x31 x21 x10      ====        or t6, s5, a0
                                                  30'd    11499    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11500    : data = 32'h    C9BF3613    ;    //    sltiu x12 x30 -869      ====        sltiu a2, t5, -869
                                                  30'd    11501    : data = 32'h    0176D613    ;    //    srli x12 x13 23      ====        srli a2, a3, 23
                                                  30'd    11502    : data = 32'h    1F3A4317    ;    //    auipc x6 127908      ====        auipc t1, 127908
                                                  30'd    11503    : data = 32'h    010A36B3    ;    //    sltu x13 x20 x16      ====        sltu a3, s4, a6
                                                  30'd    11504    : data = 32'h    414E09B3    ;    //    sub x19 x28 x20      ====        sub s3, t3, s4
                                                  30'd    11505    : data = 32'h    69A22093    ;    //    slti x1 x4 1690      ====        slti ra, tp, 1690
                                                  30'd    11506    : data = 32'h    006A5693    ;    //    srli x13 x20 6      ====        srli a3, s4, 6
                                                  30'd    11507    : data = 32'h    B84BEB93    ;    //    ori x23 x23 -1148      ====        ori s7, s7, -1148
                                                  30'd    11508    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11509    : data = 32'h    BD1F0693    ;    //    addi x13 x30 -1071      ====        addi a3, t5, -1071
                                                  30'd    11510    : data = 32'h    401DDA93    ;    //    srai x21 x27 1      ====        srai s5, s11, 1
                                                  30'd    11511    : data = 32'h    178FF493    ;    //    andi x9 x31 376      ====        andi s1, t6, 376
                                                  30'd    11512    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11513    : data = 32'h    41D5DC33    ;    //    sra x24 x11 x29      ====        sra s8, a1, t4
                                                  30'd    11514    : data = 32'h    0030E033    ;    //    or x0 x1 x3      ====        or zero, ra, gp
                                                  30'd    11515    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11516    : data = 32'h    17DECE93    ;    //    xori x29 x29 381      ====        xori t4, t4, 381
                                                  30'd    11517    : data = 32'h    9EA393B7    ;    //    lui x7 649785      ====        lui t2, 649785
                                                  30'd    11518    : data = 32'h    000A2A33    ;    //    slt x20 x20 x0      ====        slt s4, s4, zero
                                                  30'd    11519    : data = 32'h    01711FB3    ;    //    sll x31 x2 x23      ====        sll t6, sp, s7
                                                  30'd    11520    : data = 32'h    00665713    ;    //    srli x14 x12 6      ====        srli a4, a2, 6
                                                  30'd    11521    : data = 32'h    005D90B3    ;    //    sll x1 x27 x5      ====        sll ra, s11, t0
                                                  30'd    11522    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11523    : data = 32'h    006C50B3    ;    //    srl x1 x24 x6      ====        srl ra, s8, t1
                                                  30'd    11524    : data = 32'h    A8A60813    ;    //    addi x16 x12 -1398      ====        addi a6, a2, -1398
                                                  30'd    11525    : data = 32'h    005FDC33    ;    //    srl x24 x31 x5      ====        srl s8, t6, t0
                                                  30'd    11526    : data = 32'h    56846813    ;    //    ori x16 x8 1384      ====        ori a6, s0, 1384
                                                  30'd    11527    : data = 32'h    01A0FA33    ;    //    and x20 x1 x26      ====        and s4, ra, s10
                                                  30'd    11528    : data = 32'h    004CCE33    ;    //    xor x28 x25 x4      ====        xor t3, s9, tp
                                                  30'd    11529    : data = 32'h    41DD5013    ;    //    srai x0 x26 29      ====        srai zero, s10, 29
                                                  30'd    11530    : data = 32'h    40225A33    ;    //    sra x20 x4 x2      ====        sra s4, tp, sp
                                                  30'd    11531    : data = 32'h    41CD0D33    ;    //    sub x26 x26 x28      ====        sub s10, s10, t3
                                                  30'd    11532    : data = 32'h    01185413    ;    //    srli x8 x16 17      ====        srli s0, a6, 17
                                                  30'd    11533    : data = 32'h    0083EE33    ;    //    or x28 x7 x8      ====        or t3, t2, s0
                                                  30'd    11534    : data = 32'h    D9A367B7    ;    //    lui x15 891446      ====        lui a5, 891446
                                                  30'd    11535    : data = 32'h    EB223693    ;    //    sltiu x13 x4 -334      ====        sltiu a3, tp, -334
                                                  30'd    11536    : data = 32'h    D4E6E913    ;    //    ori x18 x13 -690      ====        ori s2, a3, -690
                                                  30'd    11537    : data = 32'h    E0220DB7    ;    //    lui x27 918048      ====        lui s11, 918048
                                                  30'd    11538    : data = 32'h    0105CD33    ;    //    xor x26 x11 x16      ====        xor s10, a1, a6
                                                  30'd    11539    : data = 32'h    79B70193    ;    //    addi x3 x14 1947      ====        addi gp, a4, 1947
                                                  30'd    11540    : data = 32'h    01299413    ;    //    slli x8 x19 18      ====        slli s0, s3, 18
                                                  30'd    11541    : data = 32'h    01B89E13    ;    //    slli x28 x17 27      ====        slli t3, a7, 27
                                                  30'd    11542    : data = 32'h    AFEDF313    ;    //    andi x6 x27 -1282      ====        andi t1, s11, -1282
                                                  30'd    11543    : data = 32'h    014B00B3    ;    //    add x1 x22 x20      ====        add ra, s6, s4
                                                  30'd    11544    : data = 32'h    00197A33    ;    //    and x20 x18 x1      ====        and s4, s2, ra
                                                  30'd    11545    : data = 32'h    00AF9733    ;    //    sll x14 x31 x10      ====        sll a4, t6, a0
                                                  30'd    11546    : data = 32'h    0052D8B3    ;    //    srl x17 x5 x5      ====        srl a7, t0, t0
                                                  30'd    11547    : data = 32'h    003F1FB3    ;    //    sll x31 x30 x3      ====        sll t6, t5, gp
                                                  30'd    11548    : data = 32'h    01039333    ;    //    sll x6 x7 x16      ====        sll t1, t2, a6
                                                  30'd    11549    : data = 32'h    013326B3    ;    //    slt x13 x6 x19      ====        slt a3, t1, s3
                                                  30'd    11550    : data = 32'h    00FA9EB3    ;    //    sll x29 x21 x15      ====        sll t4, s5, a5
                                                  30'd    11551    : data = 32'h    9D05CC13    ;    //    xori x24 x11 -1584      ====        xori s8, a1, -1584
                                                  30'd    11552    : data = 32'h    006BA9B3    ;    //    slt x19 x23 x6      ====        slt s3, s7, t1
                                                  30'd    11553    : data = 32'h    01AD0FB3    ;    //    add x31 x26 x26      ====        add t6, s10, s10
                                                  30'd    11554    : data = 32'h    D53773B7    ;    //    lui x7 873335      ====        lui t2, 873335
                                                  30'd    11555    : data = 32'h    009DD193    ;    //    srli x3 x27 9      ====        srli gp, s11, 9
                                                  30'd    11556    : data = 32'h    01F91AB3    ;    //    sll x21 x18 x31      ====        sll s5, s2, t6
                                                  30'd    11557    : data = 32'h    00051C13    ;    //    slli x24 x10 0      ====        slli s8, a0, 0
                                                  30'd    11558    : data = 32'h    018325B3    ;    //    slt x11 x6 x24      ====        slt a1, t1, s8
                                                  30'd    11559    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11560    : data = 32'h    4E16C313    ;    //    xori x6 x13 1249      ====        xori t1, a3, 1249
                                                  30'd    11561    : data = 32'h    01760BB3    ;    //    add x23 x12 x23      ====        add s7, a2, s7
                                                  30'd    11562    : data = 32'h    4004DA93    ;    //    srai x21 x9 0      ====        srai s5, s1, 0
                                                  30'd    11563    : data = 32'h    01BD68B3    ;    //    or x17 x26 x27      ====        or a7, s10, s11
                                                  30'd    11564    : data = 32'h    01BF4133    ;    //    xor x2 x30 x27      ====        xor sp, t5, s11
                                                  30'd    11565    : data = 32'h    01757933    ;    //    and x18 x10 x23      ====        and s2, a0, s7
                                                  30'd    11566    : data = 32'h    8E102D13    ;    //    slti x26 x0 -1823      ====        slti s10, zero, -1823
                                                  30'd    11567    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11568    : data = 32'h    0171A033    ;    //    slt x0 x3 x23      ====        slt zero, gp, s7
                                                  30'd    11569    : data = 32'h    D64C7C17    ;    //    auipc x24 877767      ====        auipc s8, 877767
                                                  30'd    11570    : data = 32'h    00789A13    ;    //    slli x20 x17 7      ====        slli s4, a7, 7
                                                  30'd    11571    : data = 32'h    0BCD1417    ;    //    auipc x8 48337      ====        auipc s0, 48337
                                                  30'd    11572    : data = 32'h    0F574B13    ;    //    xori x22 x14 245      ====        xori s6, a4, 245
                                                  30'd    11573    : data = 32'h    00B31733    ;    //    sll x14 x6 x11      ====        sll a4, t1, a1
                                                  30'd    11574    : data = 32'h    002781B3    ;    //    add x3 x15 x2      ====        add gp, a5, sp
                                                  30'd    11575    : data = 32'h    013B5193    ;    //    srli x3 x22 19      ====        srli gp, s6, 19
                                                  30'd    11576    : data = 32'h    01C77B33    ;    //    and x22 x14 x28      ====        and s6, a4, t3
                                                  30'd    11577    : data = 32'h    83CDE013    ;    //    ori x0 x27 -1988      ====        ori zero, s11, -1988
                                                  30'd    11578    : data = 32'h    FD0D3E93    ;    //    sltiu x29 x26 -48      ====        sltiu t4, s10, -48
                                                  30'd    11579    : data = 32'h    40B85193    ;    //    srai x3 x16 11      ====        srai gp, a6, 11
                                                  30'd    11580    : data = 32'h    00A5FD33    ;    //    and x26 x11 x10      ====        and s10, a1, a0
                                                  30'd    11581    : data = 32'h    010812B3    ;    //    sll x5 x16 x16      ====        sll t0, a6, a6
                                                  30'd    11582    : data = 32'h    00CC4A33    ;    //    xor x20 x24 x12      ====        xor s4, s8, a2
                                                  30'd    11583    : data = 32'h    41015B13    ;    //    srai x22 x2 16      ====        srai s6, sp, 16
                                                  30'd    11584    : data = 32'h    419C5433    ;    //    sra x8 x24 x25      ====        sra s0, s8, s9
                                                  30'd    11585    : data = 32'h    01BBA2B3    ;    //    slt x5 x23 x27      ====        slt t0, s7, s11
                                                  30'd    11586    : data = 32'h    400D8D33    ;    //    sub x26 x27 x0      ====        sub s10, s11, zero
                                                  30'd    11587    : data = 32'h    402256B3    ;    //    sra x13 x4 x2      ====        sra a3, tp, sp
                                                  30'd    11588    : data = 32'h    6E286A93    ;    //    ori x21 x16 1762      ====        ori s5, a6, 1762
                                                  30'd    11589    : data = 32'h    1E03E193    ;    //    ori x3 x7 480      ====        ori gp, t2, 480
                                                  30'd    11590    : data = 32'h    4196DD33    ;    //    sra x26 x13 x25      ====        sra s10, a3, s9
                                                  30'd    11591    : data = 32'h    01C42C33    ;    //    slt x24 x8 x28      ====        slt s8, s0, t3
                                                  30'd    11592    : data = 32'h    017F8B33    ;    //    add x22 x31 x23      ====        add s6, t6, s7
                                                  30'd    11593    : data = 32'h    01BC5193    ;    //    srli x3 x24 27      ====        srli gp, s8, 27
                                                  30'd    11594    : data = 32'h    B9107C93    ;    //    andi x25 x0 -1135      ====        andi s9, zero, -1135
                                                  30'd    11595    : data = 32'h    D3A0F413    ;    //    andi x8 x1 -710      ====        andi s0, ra, -710
                                                  30'd    11596    : data = 32'h    5A061117    ;    //    auipc x2 368737      ====        auipc sp, 368737
                                                  30'd    11597    : data = 32'h    F9244617    ;    //    auipc x12 1020484      ====        auipc a2, 1020484
                                                  30'd    11598    : data = 32'h    92780C13    ;    //    addi x24 x16 -1753      ====        addi s8, a6, -1753
                                                  30'd    11599    : data = 32'h    442B6B93    ;    //    ori x23 x22 1090      ====        ori s7, s6, 1090
                                                  30'd    11600    : data = 32'h    41C959B3    ;    //    sra x19 x18 x28      ====        sra s3, s2, t3
                                                  30'd    11601    : data = 32'h    01743FB3    ;    //    sltu x31 x8 x23      ====        sltu t6, s0, s7
                                                  30'd    11602    : data = 32'h    002AF033    ;    //    and x0 x21 x2      ====        and zero, s5, sp
                                                  30'd    11603    : data = 32'h    0078D713    ;    //    srli x14 x17 7      ====        srli a4, a7, 7
                                                  30'd    11604    : data = 32'h    CF5C0613    ;    //    addi x12 x24 -779      ====        addi a2, s8, -779
                                                  30'd    11605    : data = 32'h    01F29D33    ;    //    sll x26 x5 x31      ====        sll s10, t0, t6
                                                  30'd    11606    : data = 32'h    40148A33    ;    //    sub x20 x9 x1      ====        sub s4, s1, ra
                                                  30'd    11607    : data = 32'h    01F21A33    ;    //    sll x20 x4 x31      ====        sll s4, tp, t6
                                                  30'd    11608    : data = 32'h    01E2ACB3    ;    //    slt x25 x5 x30      ====        slt s9, t0, t5
                                                  30'd    11609    : data = 32'h    00773433    ;    //    sltu x8 x14 x7      ====        sltu s0, a4, t2
                                                  30'd    11610    : data = 32'h    D612E393    ;    //    ori x7 x5 -671      ====        ori t2, t0, -671
                                                  30'd    11611    : data = 32'h    40A80433    ;    //    sub x8 x16 x10      ====        sub s0, a6, a0
                                                  30'd    11612    : data = 32'h    00DE5913    ;    //    srli x18 x28 13      ====        srli s2, t3, 13
                                                  30'd    11613    : data = 32'h    F5F6FA13    ;    //    andi x20 x13 -161      ====        andi s4, a3, -161
                                                  30'd    11614    : data = 32'h    40185713    ;    //    srai x14 x16 1      ====        srai a4, a6, 1
                                                  30'd    11615    : data = 32'h    405304B3    ;    //    sub x9 x6 x5      ====        sub s1, t1, t0
                                                  30'd    11616    : data = 32'h    6146C293    ;    //    xori x5 x13 1556      ====        xori t0, a3, 1556
                                                  30'd    11617    : data = 32'h    00110AB3    ;    //    add x21 x2 x1      ====        add s5, sp, ra
                                                  30'd    11618    : data = 32'h    B206E993    ;    //    ori x19 x13 -1248      ====        ori s3, a3, -1248
                                                  30'd    11619    : data = 32'h    03F41D17    ;    //    auipc x26 16193      ====        auipc s10, 16193
                                                  30'd    11620    : data = 32'h    B263DDB7    ;    //    lui x27 730685      ====        lui s11, 730685
                                                  30'd    11621    : data = 32'h    00F21633    ;    //    sll x12 x4 x15      ====        sll a2, tp, a5
                                                  30'd    11622    : data = 32'h    01E8B333    ;    //    sltu x6 x17 x30      ====        sltu t1, a7, t5
                                                  30'd    11623    : data = 32'h    0177F433    ;    //    and x8 x15 x23      ====        and s0, a5, s7
                                                  30'd    11624    : data = 32'h    BFD3E593    ;    //    ori x11 x7 -1027      ====        ori a1, t2, -1027
                                                  30'd    11625    : data = 32'h    36FE0613    ;    //    addi x12 x28 879      ====        addi a2, t3, 879
                                                  30'd    11626    : data = 32'h    0042F8B3    ;    //    and x17 x5 x4      ====        and a7, t0, tp
                                                  30'd    11627    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11628    : data = 32'h    01C79B33    ;    //    sll x22 x15 x28      ====        sll s6, a5, t3
                                                  30'd    11629    : data = 32'h    40845993    ;    //    srai x19 x8 8      ====        srai s3, s0, 8
                                                  30'd    11630    : data = 32'h    010DB9B3    ;    //    sltu x19 x27 x16      ====        sltu s3, s11, a6
                                                  30'd    11631    : data = 32'h    0140D5B3    ;    //    srl x11 x1 x20      ====        srl a1, ra, s4
                                                  30'd    11632    : data = 32'h    8C223737    ;    //    lui x14 573987      ====        lui a4, 573987
                                                  30'd    11633    : data = 32'h    FFF00B93    ;    //    addi x23 x0 -1      ====        li s7, 0xffffffff #start riscv_int_numeric_corner_stream_5
                                                  30'd    11634    : data = 32'h    00000313    ;    //    addi x6 x0 0      ====        li t1, 0x0
                                                  30'd    11635    : data = 32'h    00000613    ;    //    addi x12 x0 0      ====        li a2, 0x0
                                                  30'd    11636    : data = 32'h    B10E3A37    ;    //    lui x20 725219      ====        li s4, 0xb10e33ef
                                                  30'd    11637    : data = 32'h    3EFA0A13    ;    //    addi x20 x20 1007      ====        li s4, 0xb10e33ef
                                                  30'd    11638    : data = 32'h    FFF00F93    ;    //    addi x31 x0 -1      ====        li t6, 0xffffffff
                                                  30'd    11639    : data = 32'h    FFF00B13    ;    //    addi x22 x0 -1      ====        li s6, 0xffffffff
                                                  30'd    11640    : data = 32'h    FFF00C13    ;    //    addi x24 x0 -1      ====        li s8, 0xffffffff
                                                  30'd    11641    : data = 32'h    FFF00A93    ;    //    addi x21 x0 -1      ====        li s5, 0xffffffff
                                                  30'd    11642    : data = 32'h    80000937    ;    //    lui x18 524288      ====        li s2, 0x80000000
                                                  30'd    11643    : data = 32'h    00090913    ;    //    addi x18 x18 0      ====        li s2, 0x80000000
                                                  30'd    11644    : data = 32'h    45C0F837    ;    //    lui x16 285711      ====        li a6, 0x45c0f72d
                                                  30'd    11645    : data = 32'h    72D80813    ;    //    addi x16 x16 1837      ====        li a6, 0x45c0f72d
                                                  30'd    11646    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11647    : data = 32'h    41FC0933    ;    //    sub x18 x24 x31      ====        sub s2, s8, t6
                                                  30'd    11648    : data = 32'h    3F7A0F93    ;    //    addi x31 x20 1015      ====        addi t6, s4, 1015
                                                  30'd    11649    : data = 32'h    01FA0FB3    ;    //    add x31 x20 x31      ====        add t6, s4, t6
                                                  30'd    11650    : data = 32'h    0C7B6B97    ;    //    auipc x23 51126      ====        auipc s7, 51126
                                                  30'd    11651    : data = 32'h    01230A33    ;    //    add x20 x6 x18      ====        add s4, t1, s2
                                                  30'd    11652    : data = 32'h    4990FF97    ;    //    auipc x31 301327      ====        auipc t6, 301327
                                                  30'd    11653    : data = 32'h    994B9617    ;    //    auipc x12 627897      ====        auipc a2, 627897
                                                  30'd    11654    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11655    : data = 32'h    40CC0633    ;    //    sub x12 x24 x12      ====        sub a2, s8, a2
                                                  30'd    11656    : data = 32'h    0EFF2BB7    ;    //    lui x23 61426      ====        lui s7, 61426
                                                  30'd    11657    : data = 32'h    018B8FB3    ;    //    add x31 x23 x24      ====        add t6, s7, s8
                                                  30'd    11658    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11659    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11660    : data = 32'h    016A8333    ;    //    add x6 x21 x22      ====        add t1, s5, s6
                                                  30'd    11661    : data = 32'h    10090313    ;    //    addi x6 x18 256      ====        addi t1, s2, 256
                                                  30'd    11662    : data = 32'h    BF460B93    ;    //    addi x23 x12 -1036      ====        addi s7, a2, -1036
                                                  30'd    11663    : data = 32'h    18F60313    ;    //    addi x6 x12 399      ====        addi t1, a2, 399
                                                  30'd    11664    : data = 32'h    417F8633    ;    //    sub x12 x31 x23      ====        sub a2, t6, s7
                                                  30'd    11665    : data = 32'h    3CA53A97    ;    //    auipc x21 248403      ====        auipc s5, 248403
                                                  30'd    11666    : data = 32'h    40630C33    ;    //    sub x24 x6 x6      ====        sub s8, t1, t1
                                                  30'd    11667    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11668    : data = 32'h    06BACAB7    ;    //    lui x21 27564      ====        lui s5, 27564
                                                  30'd    11669    : data = 32'h    094000EF    ;    //    jal x1 148      ====        jal storeRegisters #end riscv_int_numeric_corner_stream_5
                                                  30'd    11670    : data = 32'h    4056D5B3    ;    //    sra x11 x13 x5      ====        sra a1, a3, t0
                                                  30'd    11671    : data = 32'h    006CF4B3    ;    //    and x9 x25 x6      ====        and s1, s9, t1
                                                  30'd    11672    : data = 32'h    09CEB713    ;    //    sltiu x14 x29 156      ====        sltiu a4, t4, 156
                                                  30'd    11673    : data = 32'h    008F2CB3    ;    //    slt x25 x30 x8      ====        slt s9, t5, s0
                                                  30'd    11674    : data = 32'h    7F9E6113    ;    //    ori x2 x28 2041      ====        ori sp, t3, 2041
                                                  30'd    11675    : data = 32'h    008E1AB3    ;    //    sll x21 x28 x8      ====        sll s5, t3, s0
                                                  30'd    11676    : data = 32'h    00BDD5B3    ;    //    srl x11 x27 x11      ====        srl a1, s11, a1
                                                  30'd    11677    : data = 32'h    01812933    ;    //    slt x18 x2 x24      ====        slt s2, sp, s8
                                                  30'd    11678    : data = 32'h    41AD5393    ;    //    srai x7 x26 26      ====        srai t2, s10, 26
                                                  30'd    11679    : data = 32'h    0160F8B3    ;    //    and x17 x1 x22      ====        and a7, ra, s6
                                                  30'd    11680    : data = 32'h    40850E33    ;    //    sub x28 x10 x8      ====        sub t3, a0, s0
                                                  30'd    11681    : data = 32'h    110FE637    ;    //    lui x12 69886      ====        lui a2, 69886
                                                  30'd    11682    : data = 32'h    69722B93    ;    //    slti x23 x4 1687      ====        slti s7, tp, 1687
                                                  30'd    11683    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11684    : data = 32'h    768CEE93    ;    //    ori x29 x25 1896      ====        ori t4, s9, 1896
                                                  30'd    11685    : data = 32'h    868A4037    ;    //    lui x0 551076      ====        lui zero, 551076
                                                  30'd    11686    : data = 32'h    00EC73B3    ;    //    and x7 x24 x14      ====        and t2, s8, a4
                                                  30'd    11687    : data = 32'h    CAF5A337    ;    //    lui x6 831322      ====        lui t1, 831322
                                                  30'd    11688    : data = 32'h    00A678B3    ;    //    and x17 x12 x10      ====        and a7, a2, a0
                                                  30'd    11689    : data = 32'h    28B9B093    ;    //    sltiu x1 x19 651      ====        sltiu ra, s3, 651
                                                  30'd    11690    : data = 32'h    40D2DE93    ;    //    srai x29 x5 13      ====        srai t4, t0, 13
                                                  30'd    11691    : data = 32'h    23CEAD93    ;    //    slti x27 x29 572      ====        slti s11, t4, 572
                                                  30'd    11692    : data = 32'h    B1772E13    ;    //    slti x28 x14 -1257      ====        slti t3, a4, -1257
                                                  30'd    11693    : data = 32'h    016F7933    ;    //    and x18 x30 x22      ====        and s2, t5, s6
                                                  30'd    11694    : data = 32'h    007BD133    ;    //    srl x2 x23 x7      ====        srl sp, s7, t2
                                                  30'd    11695    : data = 32'h    01CDFDB3    ;    //    and x27 x27 x28      ====        and s11, s11, t3
                                                  30'd    11696    : data = 32'h    01E63033    ;    //    sltu x0 x12 x30      ====        sltu zero, a2, t5
                                                  30'd    11697    : data = 32'h    004C1E13    ;    //    slli x28 x24 4      ====        slli t3, s8, 4
                                                  30'd    11698    : data = 32'h    0063EAB3    ;    //    or x21 x7 x6      ====        or s5, t2, t1
                                                  30'd    11699    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11700    : data = 32'h    0000EAB3    ;    //    or x21 x1 x0      ====        or s5, ra, zero
                                                  30'd    11701    : data = 32'h    6E3AE013    ;    //    ori x0 x21 1763      ====        ori zero, s5, 1763
                                                  30'd    11702    : data = 32'h    010000EF    ;    //    jal x1 16      ====        jal storeRegisters #end riscv_int_test
                                                  30'd    11703    : data = 32'h    00000517    ;    //    auipc x10 0      ====        la x10, test_done
                                                  30'd    11704    : data = 32'h    0AC50513    ;    //    addi x10 x10 172      ====        la x10, test_done
                                                  30'd    11705    : data = 32'h    00050067    ;    //    jalr x0 x10 0      ====        jalr x0, x10, 0
                                                  30'd    11706    : data = 32'h    00010237    ;    //    lui x4 16      ====        lui x4,0x00010
                                                  30'd    11707    : data = 32'h    40020213    ;    //    addi x4 x4 1024      ====        addi x4, x4, 1024
                                                  30'd    11708    : data = 32'h    00022203    ;    //    lw x4 0(x4)      ====        lw x4, 0(x4)
                                                  30'd    11709    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11710    : data = 32'h    00122223    ;    //    sw x1 4(x4)      ====        sw x1, 4(x4)
                                                  30'd    11711    : data = 32'h    00222423    ;    //    sw x2 8(x4)      ====        sw x2, 8(x4)
                                                  30'd    11712    : data = 32'h    00322623    ;    //    sw x3 12(x4)      ====        sw x3, 12(x4)
                                                  30'd    11713    : data = 32'h    00422823    ;    //    sw x4 16(x4)      ====        sw x4, 16(x4)
                                                  30'd    11714    : data = 32'h    00522A23    ;    //    sw x5 20(x4)      ====        sw x5, 20(x4)
                                                  30'd    11715    : data = 32'h    00622C23    ;    //    sw x6 24(x4)      ====        sw x6, 24(x4)
                                                  30'd    11716    : data = 32'h    00722E23    ;    //    sw x7 28(x4)      ====        sw x7, 28(x4)
                                                  30'd    11717    : data = 32'h    02822023    ;    //    sw x8 32(x4)      ====        sw x8, 32(x4)
                                                  30'd    11718    : data = 32'h    02922223    ;    //    sw x9 36(x4)      ====        sw x9, 36(x4)
                                                  30'd    11719    : data = 32'h    02A22423    ;    //    sw x10 40(x4)      ====        sw x10, 40(x4)
                                                  30'd    11720    : data = 32'h    02B22623    ;    //    sw x11 44(x4)      ====        sw x11, 44(x4)
                                                  30'd    11721    : data = 32'h    02C22823    ;    //    sw x12 48(x4)      ====        sw x12, 48(x4)
                                                  30'd    11722    : data = 32'h    02D22A23    ;    //    sw x13 52(x4)      ====        sw x13, 52(x4)
                                                  30'd    11723    : data = 32'h    02E22C23    ;    //    sw x14 56(x4)      ====        sw x14, 56(x4)
                                                  30'd    11724    : data = 32'h    02F22E23    ;    //    sw x15 60(x4)      ====        sw x15, 60(x4)
                                                  30'd    11725    : data = 32'h    05022023    ;    //    sw x16 64(x4)      ====        sw x16, 64(x4)
                                                  30'd    11726    : data = 32'h    05122223    ;    //    sw x17 68(x4)      ====        sw x17, 68(x4)
                                                  30'd    11727    : data = 32'h    05222423    ;    //    sw x18 72(x4)      ====        sw x18, 72(x4)
                                                  30'd    11728    : data = 32'h    05322623    ;    //    sw x19 76(x4)      ====        sw x19, 76(x4)
                                                  30'd    11729    : data = 32'h    05422823    ;    //    sw x20 80(x4)      ====        sw x20, 80(x4)
                                                  30'd    11730    : data = 32'h    05522A23    ;    //    sw x21 84(x4)      ====        sw x21, 84(x4)
                                                  30'd    11731    : data = 32'h    05622C23    ;    //    sw x22 88(x4)      ====        sw x22, 88(x4)
                                                  30'd    11732    : data = 32'h    05722E23    ;    //    sw x23 92(x4)      ====        sw x23, 92(x4)
                                                  30'd    11733    : data = 32'h    07822023    ;    //    sw x24 96(x4)      ====        sw x24, 96(x4)
                                                  30'd    11734    : data = 32'h    07922223    ;    //    sw x25 100(x4)      ====        sw x25, 100(x4)
                                                  30'd    11735    : data = 32'h    07A22423    ;    //    sw x26 104(x4)      ====        sw x26, 104(x4)
                                                  30'd    11736    : data = 32'h    07B22623    ;    //    sw x27 108(x4)      ====        sw x27, 108(x4)
                                                  30'd    11737    : data = 32'h    07C22823    ;    //    sw x28 112(x4)      ====        sw x28, 112(x4)
                                                  30'd    11738    : data = 32'h    07D22A23    ;    //    sw x29 116(x4)      ====        sw x29, 116(x4)
                                                  30'd    11739    : data = 32'h    07E22C23    ;    //    sw x30 120(x4)      ====        sw x30, 120(x4)
                                                  30'd    11740    : data = 32'h    07F22E23    ;    //    sw x31 124(x4)      ====        sw x31, 124(x4)
                                                  30'd    11741    : data = 32'h    00010F37    ;    //    lui x30 16      ====        lui x30,0x00010
                                                  30'd    11742    : data = 32'h    400F0F13    ;    //    addi x30 x30 1024      ====        addi x30, x30, 1024
                                                  30'd    11743    : data = 32'h    07C20213    ;    //    addi x4 x4 124      ====        addi x4, x4, 124
                                                  30'd    11744    : data = 32'h    004F2023    ;    //    sw x4 0(x30)      ====        sw x4, 0x0(x30)
                                                  30'd    11745    : data = 32'h    00008067    ;    //    jalr x0 x1 0      ====        ret
                                                  30'd    11746    : data = 32'h    00100193    ;    //    addi x3 x0 1      ====        li gp, 1
                                                  30'd    11747    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11748    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11749    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11750    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11751    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11752    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                                                  30'd    11753    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop                                               
                                               
                                               
                                               
                                               
                                               
                                               
                                               
                                               
                                               
                               
                               
                               
                         /*      // load store test
                               
                               30'd	0	: data = 32'h	00000013	;    //	addi x0 x0 0	  ====    	nop
                               30'd    1    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                               30'd    2    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                               30'd    3    : data = 32'h    000000B7    ;    //    lui x1 0      ====        lui x1, 0x00000
                               30'd    4    : data = 32'h    40008093    ;    //    addi x1 x1 1024      ====        addi x1, x1, 1024
                               30'd    5    : data = 32'h    22222137    ;    //    lui x2 139810      ====        lui x2, 0x22222
                               30'd    6    : data = 32'h    0020A223    ;    //    sw x2 4(x1)      ====        sw x2, 4(x1)
                               30'd    7    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    8    : data = 32'h    333331B7    ;    //    lui x3 209715      ====        lui x3, 0x33333
                               30'd    9    : data = 32'h    0030A223    ;    //    sw x3 4(x1)      ====        sw x3, 4(x1)
                               30'd    10    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    11    : data = 32'h    44444237    ;    //    lui x4 279620      ====        lui x4, 0x44444
                               30'd    12    : data = 32'h    0040A223    ;    //    sw x4 4(x1)      ====        sw x4, 4(x1)
                               30'd    13    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    14    : data = 32'h    555552B7    ;    //    lui x5 349525      ====        lui x5, 0x55555
                               30'd    15    : data = 32'h    0050A223    ;    //    sw x5 4(x1)      ====        sw x5, 4(x1)
                               30'd    16    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    17    : data = 32'h    66666337    ;    //    lui x6 419430      ====        lui x6, 0x66666
                               30'd    18    : data = 32'h    0060A223    ;    //    sw x6 4(x1)      ====        sw x6, 4(x1)
                               30'd    19    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    20    : data = 32'h    777773B7    ;    //    lui x7 489335      ====        lui x7, 0x77777
                               30'd    21    : data = 32'h    0070A223    ;    //    sw x7 4(x1)      ====        sw x7, 4(x1)
                               30'd    22    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    23    : data = 32'h    88888437    ;    //    lui x8 559240      ====        lui x8, 0x88888
                               30'd    24    : data = 32'h    0080A223    ;    //    sw x8 4(x1)      ====        sw x8, 4(x1)
                               30'd    25    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    26    : data = 32'h    999904B7    ;    //    lui x9 629136      ====        lui x9, 0x99990
                               30'd    27    : data = 32'h    0090A223    ;    //    sw x9 4(x1)      ====        sw x9, 4(x1)
                               30'd    28    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    29    : data = 32'h    000000B7    ;    //    lui x1 0      ====        lui x1, 0x00000
                               30'd    30    : data = 32'h    40008093    ;    //    addi x1 x1 1024      ====        addi x1, x1, 1024
                               30'd    31    : data = 32'h    0040A503    ;    //    lw x10 4(x1)      ====        lw x10, 4(x1)
                               30'd    32    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    33    : data = 32'h    0040A583    ;    //    lw x11 4(x1)      ====        lw x11, 4(x1)
                               30'd    34    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    35    : data = 32'h    0040A603    ;    //    lw x12 4(x1)      ====        lw x12, 4(x1)
                               30'd    36    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    37    : data = 32'h    0040A683    ;    //    lw x13 4(x1)      ====        lw x13, 4(x1)
                               30'd    38    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    39    : data = 32'h    0040A703    ;    //    lw x14 4(x1)      ====        lw x14, 4(x1)
                               30'd    40    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    41    : data = 32'h    0040A783    ;    //    lw x15 4(x1)      ====        lw x15, 4(x1)
                               30'd    42    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    43    : data = 32'h    0040A803    ;    //    lw x16 4(x1)      ====        lw x16, 4(x1)
                               30'd    44    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    45    : data = 32'h    0040A883    ;    //    lw x17 4(x1)      ====        lw x17, 4(x1)
                               30'd    46    : data = 32'h    00408093    ;    //    addi x1 x1 4      ====        addi x1, x1, 4
                               30'd    47    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                               30'd    48    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                               30'd    49    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop
                               
                               
                              
                               */
                               
                               
                               
                               
                               
                               
	
	/*	                       
            30'd	0	: data = 32'h	FFF00813	;    //	addi x16 x0 -1	  ====    	li a6, 0xffffffff	
            30'd    1    : data = 32'h    00000513    ;    //    addi x10 x0 0      ====        li a0, 0x0    
            30'd    2    : data = 32'h    FFF00293    ;    //    addi x5 x0 -1      ====        li t0, 0xffffffff    
            30'd    3    : data = 32'h    FFF00693    ;    //    addi x13 x0 -1      ====        li a3, 0xffffffff    
            30'd    4    : data = 32'h    3CE65C37    ;    //    lui x24 249445      ====        li s8, 0x3ce64b2f    
            30'd    5    : data = 32'h    B2FC0C13    ;    //    addi x24 x24 -1233      ====        li s8, 0x3ce64b2f    
            30'd    6    : data = 32'h    00000193    ;    //    addi x3 x0 0      ====        li gp, 0x0    
            30'd    7    : data = 32'h    997F4637    ;    //    lui x12 628724      ====        li a2, 0x997f3afc    
            30'd    8    : data = 32'h    AFC60613    ;    //    addi x12 x12 -1284      ====        li a2, 0x997f3afc    
            30'd    9    : data = 32'h    00000393    ;    //    addi x7 x0 0      ====        li t2, 0x0    
            30'd    10    : data = 32'h    FFF00E13    ;    //    addi x28 x0 -1      ====        li t3, 0xffffffff    
            30'd    11    : data = 32'h    F71B26B7    ;    //    lui x13 1012146      ====        lui a3, 1012146    
            30'd    12    : data = 32'h    07660813    ;    //    addi x16 x12 118      ====        addi a6, a2, 118    
            30'd    13    : data = 32'h    CF280613    ;    //    addi x12 x16 -782      ====        addi a2, a6, -782    
            30'd    14    : data = 32'h    CE2BCE17    ;    //    auipc x28 844476      ====        auipc t3, 844476    
            30'd    15    : data = 32'h    51668E13    ;    //    addi x28 x13 1302      ====        addi t3, a3, 1302    
            30'd    16    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop    
            30'd    17    : data = 32'h    00000013    ;    //    addi x0 x0 0      ====        nop    

			
			
		
			30'h00000000: data = 32'hFFF00813; 
			30'h00000001: data = 32'h00000513; 
			30'h00000002: data = 32'h10110111; 
			30'h00000003: data = 32'h10011111; 
			30'h00000004: data = 32'h11001101; 
			30'h00000005: data = 32'h11011011; 
			30'h00000006: data = 32'h11111011; 
			30'h00000007: data = 32'h00001111; 
			30'h00000008: data = 32'h11111111; 
			30'h00000009: data = 32'h11011111; 
			*/
			30'd    12000    : $finish;
			 	 default: data = 32'h00000013; 
 		endcase

	assign irdata_o = ird_i ? data : 32'h0;
endmodule